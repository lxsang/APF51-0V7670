library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity imx_in is
  port (
    reset: in std_logic;
	clk:in std_logic;
    start: in std_logic;
	da  : out std_logic_vector(15 downto 0);
    --ready  : out std_logic;
    adv    : out std_logic;
    cs     : out std_logic;
    rw     : out std_logic;
    finish : in std_logic
  ) ;
end entity imx_in;

architecture arch of imx_in is
  type ram_type is array (0 to 2**14-1) of std_logic_vector(15 downto 0) ;
  
	signal ram:ram_type  := (

      X"D5D8",X"D4D4",X"D5D5",X"D2D2",X"DFD5",X"D3DE",X"CACC",X"D0CB",
      X"E0D5",X"DEE5",X"D0D4",X"CBCE",X"D9D2",X"E1E1",X"CDD7",X"D3CE",
      X"999E",X"FFDC",X"FFFF",X"FFFE",X"FDFD",X"FDFE",X"F9FD",X"FCFB",
      X"FCF9",X"FBFB",X"FBF9",X"FBF9",X"FCFC",X"F8F9",X"DEED",X"F7E3",
      X"FAFF",X"F8F9",X"FBFB",X"FCF9",X"F7F9",X"FBF9",X"FBFB",X"FCFB",
      X"FCFE",X"FFFF",X"B9F2",X"999A",X"9099",X"8F8D",X"8D8F",X"978F",
      X"D2C5",X"CECE",X"D5D8",X"D4D4",X"D5D5",X"D2D2",X"DFD5",X"D3DE",
      X"CACC",X"D0CB",X"E0D5",X"DEE5",X"D0D4",X"CBCE",X"D9D2",X"E1E1",
      X"D6DA",X"CDD2",X"CDCD",X"CECE",X"DAD2",X"CFD7",X"CDCC",X"CECE",
      X"D7CF",X"D5DA",X"CFCD",X"CFCF",X"D3CF",X"DBD9",X"D0D6",X"8ABA",
      X"FEBE",X"FFFF",X"FBFD",X"FAFD",X"FAFC",X"FDFB",X"FAFA",X"FEFC",
      X"FDFD",X"F9FA",X"FBF9",X"FCFB",X"F9F9",X"FAFB",X"EDF9",X"CFDA",
      X"FFE5",X"FBFE",X"FBF9",X"F9FC",X"F9FB",X"FCF9",X"F9FB",X"FAF9",
      X"FCFA",X"FEFD",X"FFFF",X"ABE4",X"9191",X"8E8B",X"8D90",X"928F",
      X"A490",X"CFC8",X"D6DA",X"CDD2",X"CDCD",X"CECE",X"DAD2",X"CFD7",
      X"CDCC",X"CECE",X"D7CF",X"D5DA",X"CFCD",X"CFCF",X"D3CF",X"DBD9",
      X"D9DE",X"CBD2",X"C9C8",X"CECB",X"D6D3",X"CED4",X"D0CD",X"CECD",
      X"D3CD",X"CFD4",X"CDCC",X"CECE",X"D2CE",X"D9D6",X"86C9",X"E28C",
      X"FFFF",X"FAFE",X"FBFB",X"FCFC",X"FCFC",X"FDFA",X"FCFA",X"FAFC",
      X"FDFC",X"FAFD",X"F9F9",X"F9FC",X"FBFB",X"FCFC",X"FEFD",X"E8FC",
      X"D3C9",X"FFF8",X"F9FC",X"F9F9",X"FDFA",X"FCFD",X"FCFC",X"FAFD",
      X"FAFA",X"FEFD",X"FEFE",X"FCFF",X"95C2",X"8B8E",X"8E8D",X"938E",
      X"9090",X"B791",X"D9DE",X"CBD2",X"C9C8",X"CECB",X"D6D3",X"CED4",
      X"D0CD",X"CECD",X"D3CD",X"CFD4",X"CDCC",X"CECE",X"D2CE",X"D9D6",
      X"DBDF",X"CFD6",X"CCCC",X"D1CE",X"DAD7",X"D1D6",X"D1D2",X"CED0",
      X"D7D5",X"D5D8",X"CDD0",X"C7CB",X"D8D1",X"CCDF",X"A766",X"FFF9",
      X"FDFE",X"FBFB",X"FBF9",X"FAFA",X"FBFA",X"FDFA",X"FCFC",X"FCFA",
      X"FDFA",X"FCFA",X"FBF9",X"F9F9",X"F9F9",X"FBFB",X"FBFB",X"FFFB",
      X"C1F4",X"EABC",X"FEFF",X"FDFD",X"FAFD",X"FAFA",X"FDFD",X"FDFD",
      X"FAFA",X"FDFD",X"FBFC",X"FEFA",X"DAFF",X"968F",X"8C8A",X"928E",
      X"9394",X"8A8E",X"DBBB",X"CFD6",X"CCCC",X"D1CE",X"DAD7",X"D1D6",
      X"D1D2",X"CED0",X"D7D5",X"D5D8",X"CDD0",X"C7CB",X"D8D1",X"DDDF",
      X"DBDB",X"D5D9",X"D1D2",X"D6D4",X"DFD9",X"D8DE",X"D4D6",X"D8D4",
      X"DEDF",X"DCDE",X"D2D8",X"C9CD",X"DFD8",X"65C5",X"FFC7",X"FEFF",
      X"FBFD",X"FBFC",X"FDFB",X"F9FF",X"FAFD",X"FAFC",X"FBFC",X"FCFC",
      X"F9FC",X"FBFB",X"FBFB",X"FBFB",X"F9FB",X"F9F9",X"FBFB",X"FCF9",
      X"F8FF",X"B5CC",X"FFDA",X"FEFF",X"FBFC",X"FEFA",X"FCFD",X"FAFC",
      X"F9FC",X"F9FA",X"FAF9",X"F9FA",X"FFFD",X"83E4",X"9090",X"9593",
      X"9696",X"8F92",X"AD93",X"D5D9",X"D1D2",X"D6D4",X"DFD9",X"D8DE",
      X"D4D6",X"D8D4",X"DEDF",X"DCDE",X"D2D8",X"C9CD",X"DFD8",X"E2E4",
      X"D9D7",X"D8D9",X"D3D6",X"D7D5",X"E0D9",X"DDE1",X"D8DA",X"DFD8",
      X"DFE2",X"DFDE",X"D8DD",X"D6D5",X"9FDF",X"DC78",X"FFFF",X"FCFD",
      X"F9FC",X"FBFB",X"FEFE",X"E9E0",X"FBFD",X"FBF9",X"FCFC",X"FBF9",
      X"FBFA",X"FBFA",X"FBF9",X"FCFB",X"FBFC",X"FBFB",X"FBFB",X"FBFB",
      X"FEFA",X"E3FF",X"C6B2",X"FFFD",X"F9FA",X"FCFC",X"FBFC",X"FBF8",
      X"F9FC",X"F9FA",X"F9FC",X"F9F9",X"FEFA",X"E2FF",X"9975",X"9797",
      X"9694",X"9697",X"9390",X"D8BE",X"D3D6",X"D7D5",X"E0D9",X"DDE1",
      X"D8DA",X"DFD8",X"DFE2",X"DFDE",X"D8DD",X"D6D5",X"E0DF",X"E4E4",
      X"D9D7",X"D8D9",X"D2D4",X"D9D5",X"DFD9",X"DDE0",X"D8DB",X"DFD8",
      X"DEE2",X"DFDC",X"D8DD",X"DAD8",X"8C97",X"FFF0",X"FDFF",X"FDFC",
      X"FBFA",X"FFF9",X"D3FF",X"F3C5",X"FBFD",X"F9F9",X"F9FB",X"F9FB",
      X"F9FB",X"FBFB",X"FBFB",X"FCF9",X"F9FC",X"F9F9",X"F9FB",X"F9FB",
      X"FCFB",X"FFFC",X"B0EB",X"FCBF",X"F8FF",X"FAFA",X"FCFB",X"FCFA",
      X"FAFC",X"F9F9",X"FBF9",X"F8F9",X"FAF9",X"FFFE",X"77C3",X"999A",
      X"9593",X"9896",X"9390",X"D699",X"D2D4",X"D9D5",X"DFD9",X"DDE0",
      X"D8DB",X"DFD8",X"DEE2",X"DFDC",X"D8DD",X"DBD8",X"E1DF",X"E3E3",
      X"DBD9",X"D8DB",X"D2D4",X"D9D7",X"DFDC",X"DCDF",X"D7DA",X"D9D6",
      X"DDE1",X"DFDD",X"D7DD",X"8BD1",X"FEA2",X"FFFF",X"FCFE",X"FAFC",
      X"FBFA",X"FFFB",X"B6DB",X"FEEE",X"F8F8",X"F9F9",X"FBFB",X"F9FB",
      X"F8F7",X"F9F8",X"FBFB",X"FBFB",X"FCFB",X"FAFA",X"F9FB",X"FBF9",
      X"FCFB",X"FBF9",X"F1FF",X"BEB6",X"FFF7",X"F9FB",X"FDFB",X"FBFC",
      X"FBF9",X"FAF9",X"F9F9",X"F9F7",X"F8F8",X"FFF8",X"94FF",X"9791",
      X"9595",X"9294",X"9391",X"B195",X"D2D4",X"D9D7",X"DFDC",X"DCDF",
      X"D7DA",X"D9D6",X"DDE1",X"DFDD",X"D7DD",X"D7D4",X"E2DC",X"E3E6",
      X"DCDD",X"D3D8",X"CCCD",X"D5D0",X"E0DC",X"D7DE",X"CCD1",X"D4CE",
      X"DCDC",X"DEDE",X"D0DA",X"A789",X"FFFF",X"FBFE",X"F9F9",X"F9FA",
      X"FAFC",X"E5FF",X"E1AF",X"FBFF",X"FAF8",X"FAF8",X"F9F9",X"F9F9",
      X"F9FB",X"F9F8",X"FBF9",X"FAFA",X"FCFA",X"FBFC",X"FBFB",X"F9F9",
      X"FBFB",X"F7F9",X"FFFB",X"AFF2",X"F8B9",X"FAFF",X"FBF9",X"FBFB",
      X"F7F9",X"F9F9",X"F8FA",X"F8F7",X"F7F8",X"FBF7",X"DEFF",X"9984",
      X"9797",X"8F94",X"9694",X"9294",X"CCC5",X"D5D0",X"E0DC",X"D7DE",
      X"CCD1",X"D4CE",X"DCDC",X"DEDE",X"D3DA",X"CFD0",X"DED6",X"E0E2",
      X"D9DD",X"CAD2",X"C4C6",X"C9C7",X"DFD8",X"D1DC",X"CACB",X"CECA",
      X"DCD5",X"D8DE",X"87CE",X"FFAE",X"FEFF",X"FAFB",X"FBF9",X"F9FA",
      X"FFFD",X"B2F3",X"FFD8",X"FAFC",X"FAFA",X"F9FA",X"FBF9",X"FBF9",
      X"F9FB",X"F9FA",X"F9F9",X"F9F9",X"F9F9",X"F9F9",X"F9F9",X"F8F8",
      X"F8F9",X"F9FA",X"F9F9",X"ECFF",X"C1B4",X"FEFC",X"F9F9",X"F9F9",
      X"FAF8",X"FBFA",X"F8F9",X"F8F7",X"F7F8",X"F7F9",X"FFFC",X"94B0",
      X"9294",X"9092",X"9394",X"8C90",X"C49F",X"C9C7",X"DFD8",X"D1DC",
      X"CACB",X"CECA",X"DCD5",X"D8DE",X"CFD1",X"CCCD",X"D7CF",X"D8D9",
      X"D5DA",X"C8CF",X"C5C5",X"C9C8",X"DED5",X"D1DD",X"CDCC",X"D0CE",
      X"D9CF",X"D0DB",X"A987",X"FFFF",X"FAFC",X"FBF9",X"FAFB",X"FAFC",
      X"FDFE",X"BFB5",X"FEFF",X"FBFA",X"FBFC",X"FBFB",X"FBF9",X"F9FB",
      X"F8F9",X"F9F9",X"F8F9",X"F9FA",X"F9FA",X"F9F7",X"F9F9",X"F8F8",
      X"F7F8",X"F6F6",X"F6F7",X"FDF7",X"B5F0",X"FBC7",X"F7FD",X"F7F7",
      X"FBF7",X"F9FB",X"F8F9",X"F8F8",X"F6F7",X"F9F8",X"FFF9",X"84EA",
      X"9199",X"928F",X"9093",X"8B8E",X"BB8A",X"C9C8",X"DED5",X"D1DD",
      X"CDCC",X"D0CE",X"D9CF",X"D4DB",X"CCCB",X"D0CE",X"D6CE",X"D8DA",
      X"D6D8",X"CDD2",X"CAC9",X"D0CD",X"E0D8",X"D6DF",X"CFD0",X"D2CF",
      X"D9D3",X"7FD6",X"FFB4",X"FAFF",X"FCF9",X"FCFA",X"FAFC",X"FCFC",
      X"CDFF",X"F4A6",X"FCFF",X"FBFA",X"FDFB",X"FBFB",X"F9F9",X"F8FA",
      X"F9F7",X"F7F9",X"FAF7",X"F8F7",X"F7F8",X"F7F8",X"F6F7",X"F6F7",
      X"F7F7",X"F7F6",X"F7F6",X"F9F7",X"EFFE",X"C6B4",X"FCFE",X"F7F9",
      X"F9F7",X"FAFB",X"F7F7",X"F7F7",X"F9F7",X"F6F6",X"FBF7",X"ABFF",
      X"9292",X"8D8F",X"9292",X"8F91",X"9E8D",X"D0CD",X"E0D8",X"D6DF",
      X"CFD0",X"D2CF",X"D9D3",X"D6DC",X"CDCE",X"D0CF",X"DCD2",X"DBE0",
      X"D9D8",X"D5DA",X"CCCF",X"D5D0",X"E0DE",X"DCDF",X"CFD8",X"D2CD",
      X"DDDE",X"A877",X"FFFF",X"FBFD",X"FCFB",X"F9FC",X"FCF9",X"FFFC",
      X"A0E9",X"FFDF",X"FBFC",X"FBFA",X"F9FA",X"F8FA",X"F8F7",X"F9FA",
      X"F9F9",X"F8F7",X"FAF8",X"FCFC",X"F8FB",X"F8F8",X"F7F6",X"F7F7",
      X"F8F6",X"F7F8",X"F8F8",X"F5F7",X"FEF9",X"AFEA",X"FFCF",X"F8FA",
      X"F7F7",X"F8F8",X"F7F7",X"F7F7",X"F6F7",X"F7F6",X"F6F6",X"E9FF",
      X"9D87",X"9294",X"9392",X"9495",X"8D90",X"D5C3",X"E0DE",X"DCDF",
      X"CFD8",X"D2CD",X"DDDE",X"DDDE",X"D1D9",X"D3CF",X"DED9",X"DBDE",
      X"DDD9",X"DDE1",X"D5D7",X"DED9",X"E0DF",X"E1DF",X"D6DF",X"DBD4",
      X"8FE1",X"FF95",X"FCFF",X"FBFB",X"FCFB",X"FAFC",X"FBFA",X"FBFE",
      X"BDB3",X"FEFF",X"F9F9",X"F8F8",X"F7F7",X"F7F7",X"F6F7",X"F7F6",
      X"FAF8",X"F7F8",X"FBF7",X"EEF6",X"FAFB",X"F7F7",X"F7F7",X"FAFB",
      X"F6F7",X"F7F7",X"F6F7",X"F4F6",X"F8F7",X"DEFF",X"DAA4",X"F6FE",
      X"F7F7",X"F7F7",X"F7F8",X"F7F8",X"F8F6",X"F5F5",X"F5F5",X"FFFB",
      X"90B5",X"9698",X"9692",X"979A",X"9295",X"DEA5",X"E0DF",X"E1DF",
      X"D6DF",X"DBD4",X"DDE1",X"E2DE",X"D9E0",X"D9D5",X"E0DF",X"DCDD",
      X"DDDA",X"DFE0",X"DAD9",X"E3DE",X"E0DE",X"E1E0",X"DBE0",X"E1DA",
      X"76B9",X"FFF0",X"F9FB",X"FBFB",X"F9F9",X"F9FC",X"FBF9",X"D5FF",
      X"F2A5",X"FAFF",X"F7F9",X"F9F9",X"F9F8",X"F8FA",X"F8FB",X"F7F7",
      X"F8F8",X"F7F7",X"F9F6",X"C6E7",X"FBF5",X"F8F7",X"F9F9",X"F6F7",
      X"F6FA",X"F7F6",X"F6F8",X"F8F7",X"F5F9",X"FFF8",X"A0CD",X"FBEA",
      X"F6F6",X"F7F7",X"F7F8",X"F6F1",X"F4F9",X"F5F4",X"F5F5",X"FFF6",
      X"8BEE",X"979C",X"9391",X"9896",X"9494",X"D396",X"E0DE",X"E1E0",
      X"DBE0",X"E1DA",X"DEDF",X"E1DF",X"DCE0",X"DAD9",X"E1E0",X"E0DF",
      X"DDDC",X"DADD",X"D6D6",X"DCD8",X"E3DF",X"DEE2",X"D8DA",X"D5D6",
      X"E383",X"FDFF",X"FBF9",X"F8F9",X"FBF7",X"F9FB",X"FFF9",X"A7F4",
      X"FFD0",X"F9F9",X"F7F7",X"F7F7",X"F6F8",X"FBF9",X"F2FA",X"F7F8",
      X"F8F8",X"F8F8",X"FBF4",X"BCDF",X"FBF7",X"F8F8",X"F7FB",X"E7CC",
      X"F8FD",X"F6F7",X"F9F9",X"F8F7",X"F6F9",X"FCF6",X"BCFD",X"F4B3",
      X"F5FA",X"F8F7",X"F6FA",X"ECDA",X"F5F8",X"F4F4",X"F5F4",X"FAF3",
      X"B7FF",X"948C",X"9391",X"9394",X"9091",X"A48F",X"E3DF",X"DEE2",
      X"D8DA",X"DAD6",X"E3E0",X"E0E5",X"D8DC",X"D5D6",X"DFD8",X"E0E1",
      X"DADC",X"D6D9",X"CED1",X"D4D0",X"E1D9",X"DFE4",X"D0D7",X"9CCE",
      X"FFDA",X"FBFD",X"FAFB",X"F7FA",X"FAF8",X"F8F9",X"FFF9",X"A9C7",
      X"FCF8",X"F7F7",X"F7F7",X"F8F7",X"F6F7",X"FEF9",X"DCDC",X"F9FB",
      X"F7F7",X"F8F9",X"FDF7",X"C5DE",X"FBFA",X"F7F7",X"FAFC",X"D09F",
      X"F5FF",X"F7F6",X"F4F0",X"F6FA",X"F5F6",X"F8F6",X"F3FE",X"B8AF",
      X"FAF7",X"F6F5",X"FBF9",X"D1D2",X"F6F9",X"F3F4",X"F4F3",X"F4F2",
      X"EAFE",X"9381",X"9395",X"9294",X"8E8F",X"908E",X"E1CB",X"DFE4",
      X"D0D7",X"D4CE",X"DEDC",X"E1E3",X"D1D7",X"CBD0",X"D9D7",X"E1E1",
      X"D7D9",X"D2D4",X"CBCE",X"D1CD",X"DED9",X"D5DB",X"CED2",X"CAA7",
      X"FDFF",X"FCFC",X"FAFA",X"F9F8",X"F8F7",X"F9F8",X"EBFF",X"DB9C",
      X"F7FF",X"F6F7",X"FAF9",X"F7F9",X"F6F7",X"EDFB",X"E4BB",X"F5FD",
      X"F7F5",X"F8F7",X"FEFA",X"BADB",X"FBF9",X"F6F7",X"FEFC",X"C18D",
      X"F4FF",X"F9F6",X"D4E0",X"F9F7",X"F5F3",X"F7F7",X"FEF7",X"99E9",
      X"FEBC",X"F4F9",X"FDF6",X"B8E1",X"F7EE",X"F3F3",X"F2F2",X"F2F2",
      X"FFF9",X"86B5",X"9393",X"9291",X"8C8F",X"8F8E",X"DEA3",X"D5DB",
      X"CED2",X"CECD",X"D9D7",X"D9DD",X"CDD2",X"CBCF",X"D3CF",X"DADB",
      X"D6DA",X"D0D2",X"CBCC",X"D0CC",X"D8D5",X"CFD5",X"A8CD",X"FFB4",
      X"F7FE",X"F9F9",X"FBFB",X"F1EF",X"F8FA",X"FCF8",X"AEFF",X"FFB1",
      X"F8FE",X"F8F6",X"F9FA",X"F7F8",X"F8F7",X"CEFD",X"FEC0",X"F6FB",
      X"F7F5",X"F7F7",X"FFFA",X"AFD0",X"FBFB",X"F5F6",X"FCFB",X"C28D",
      X"F6FF",X"FCF5",X"C0EF",X"FBDA",X"F2F5",X"F7F5",X"F6F5",X"D6FF",
      X"D893",X"F6FF",X"F9F5",X"B7F1",X"FBDB",X"F4F5",X"F2F2",X"F2F1",
      X"FCF5",X"92F7",X"9298",X"9192",X"8D8E",X"8F8E",X"C193",X"CFD5",
      X"CDCD",X"CDCC",X"D4CF",X"D5D9",X"CDCF",X"CDD0",X"D1CB",X"D8D8",
      X"D7DC",X"CFD3",X"C9CB",X"CFCB",X"DBD2",X"D4DB",X"94AD",X"FFFD",
      X"F7F8",X"F7F9",X"FCFB",X"DBC6",X"F8FC",X"FFFA",X"9FDC",X"FFEB",
      X"F3EC",X"F7FB",X"F7F8",X"F7F8",X"FBF7",X"BDFB",X"FED9",X"F7F9",
      X"F8F7",X"F7F7",X"FFF9",X"B1CC",X"F9FC",X"F5F4",X"FDFB",X"C590",
      X"F7FF",X"F6F6",X"DAFC",X"EEBD",X"F4F9",X"F5F3",X"F4F5",X"FCF7",
      X"9DC0",X"FEEC",X"F6F3",X"C4FB",X"F9C0",X"F4F4",X"F1F1",X"EFF0",
      X"F3F0",X"CBFE",X"9393",X"8F91",X"8C8D",X"8E8C",X"A490",X"D4DB",
      X"CBCE",X"CECC",X"D6D0",X"D8DC",X"CFD1",X"CCCE",X"D5CE",X"DADC",
      X"D6DA",X"D0D3",X"CCCE",X"D4CF",X"E3DC",X"CFE0",X"ED80",X"FBFF",
      X"F7F9",X"F8F8",X"F3FC",X"DEB1",X"F7FC",X"F8FD",X"CBAF",X"F1FF",
      X"F5D5",X"F7FA",X"F9F7",X"F7F8",X"FFF9",X"BBE4",X"FBF1",X"F7F9",
      X"F7F7",X"F7F7",X"FEF6",X"B6CE",X"F8FC",X"F5F4",X"FEFD",X"BF93",
      X"F6FF",X"F4F5",X"F5F5",X"CCBD",X"F3F9",X"F4F2",X"F4F3",X"F8F4",
      X"A1EF",X"FEBB",X"F3F6",X"DAFA",X"EDA9",X"F2F6",X"F1F1",X"EFF0",
      X"F1F0",X"F3F9",X"9696",X"8E90",X"8B8D",X"908D",X"9996",X"D8C2",
      X"D1D4",X"D1CF",X"E0D9",X"DEE2",X"D1D6",X"CCCE",X"DBD4",X"DFE0",
      X"D9DC",X"D8D8",X"D5D5",X"DFDA",X"E2E5",X"68DC",X"FFC9",X"F9FB",
      X"F7F9",X"F7F6",X"E5FD",X"EEAE",X"F7FC",X"DBFF",X"F0A8",X"DBFF",
      X"F9E2",X"F9F8",X"F8F7",X"F8F8",X"FDF9",X"CEC7",X"F4FA",X"F7F7",
      X"F6F6",X"F6F7",X"FEF7",X"B0C6",X"F9FE",X"F4F5",X"FFFD",X"B88E",
      X"F6FF",X"F0F3",X"F9F1",X"B4D6",X"F6EA",X"F2F1",X"F1F2",X"F3F1",
      X"DDFB",X"DA9A",X"F1FD",X"EDF7",X"DAA1",X"F2F7",X"F2F1",X"F0F0",
      X"F0F0",X"FBF2",X"7CC9",X"9395",X"9191",X"9693",X"979B",X"D496",
      X"D9DB",X"D9D8",X"E2E0",X"DFE3",X"D7DC",X"D8D5",X"DFD9",X"E2E2",
      X"DDDD",X"DCDE",X"D9DA",X"E5DE",X"E0E4",X"96AB",X"FDFF",X"F8F7",
      X"F8F8",X"F7F6",X"D5FD",X"FCB6",X"FBF8",X"BCFB",X"FFCF",X"CAED",
      X"F9F4",X"F8F8",X"F6F8",X"F7F7",X"F2FA",X"E5B6",X"F2FA",X"F6F6",
      X"F7F5",X"F6F6",X"FFFA",X"B5B7",X"F7FF",X"F4F6",X"FEF9",X"B387",
      X"F5FF",X"EEF1",X"F4EF",X"BBED",X"F8D1",X"F0F0",X"F0F0",X"F1EE",
      X"FBF4",X"9AB6",X"FAED",X"F7F6",X"C2AD",X"F1F9",X"F1F1",X"F0F1",
      X"EFF0",X"F3EF",X"9EF6",X"968B",X"9394",X"9B96",X"9699",X"AA92",
      X"DCDD",X"DDD9",X"E0DF",X"E0DF",X"DBE0",X"DED9",X"E2DF",X"E1E0",
      X"DBDA",X"DBDD",X"D3D6",X"DFD7",X"DCE3",X"E975",X"F7FF",X"F7F7",
      X"F8F8",X"F8F6",X"C3FF",X"FFC1",X"FFF7",X"ADD8",X"FFF3",X"D0D0",
      X"F9FE",X"F8F8",X"F6F8",X"F6F7",X"DEFD",X"F2B4",X"F2F3",X"F5F5",
      X"F3F3",X"F5F5",X"FBF7",X"C4B3",X"F5FE",X"F5F5",X"FBFB",X"B884",
      X"F3FF",X"E9F1",X"EFE6",X"D3F8",X"F1B5",X"F0F7",X"F0EF",X"EFEF",
      X"F8EE",X"95E8",X"FBBC",X"FAF3",X"B7C7",X"F0F5",X"EEEE",X"EFEF",
      X"EDF0",X"EEEC",X"E7F5",X"9A8F",X"8F92",X"9693",X"979A",X"9796",
      X"D5C0",X"D8D2",X"E0E1",X"E3DF",X"DCE4",X"DCD6",X"E3E3",X"DCDD",
      X"D9DE",X"D3D6",X"CCCD",X"D8D2",X"BEDE",X"FF94",X"F9FB",X"F9F7",
      X"F8F8",X"FCF6",X"ADFC",X"FFCB",X"F9FB",X"C9AD",X"EDFF",X"E7BC",
      X"F4FC",X"F8F7",X"F4F8",X"F7F5",X"CCFC",X"F2BE",X"EEDD",X"F4F5",
      X"F2F3",X"F0F1",X"F6F2",X"CFB1",X"F5FE",X"F4F4",X"F8FC",X"C88F",
      X"F4FE",X"EFF1",X"E3E1",X"E8F5",X"DFA9",X"F0FD",X"F0EF",X"EFF1",
      X"EFEF",X"D0F9",X"E495",X"F9F9",X"ABD9",X"F3E9",X"EBEC",X"EDEC",
      X"EFEE",X"EAEC",X"F9EC",X"91D8",X"8C91",X"938F",X"9A96",X"9399",
      X"C490",X"D2CE",X"DDD7",X"DFE1",X"D6DA",X"CFD1",X"DAD8",X"DFE0",
      X"D6D9",X"CED2",X"C5C8",X"D1CB",X"8BDB",X"FFC2",X"F9F8",X"F9F7",
      X"F7F9",X"FCF7",X"A5F4",X"FDD6",X"D5FC",X"F0A6",X"CBFF",X"FBC9",
      X"F4F6",X"F5F6",X"F4F4",X"F6F6",X"C1F8",X"DFD9",X"F3B7",X"F3F9",
      X"F1F3",X"EFF0",X"F2F6",X"D2A7",X"F4FF",X"F2F2",X"F2F9",X"D493",
      X"F1FC",X"F1EF",X"D9EB",X"F8E3",X"BBC1",X"F5F7",X"F2F0",X"EFF2",
      X"EDED",X"F2F2",X"B5A1",X"F8F7",X"A2E7",X"F6DD",X"ECEB",X"EDEC",
      X"EEED",X"EBEB",X"D8EB",X"CFEB",X"8A94",X"8F8C",X"9795",X"9095",
      X"958D",X"C8C5",X"D9D3",X"DADD",X"CDD2",X"CCCB",X"D3CE",X"DBDB",
      X"D6DA",X"CBD0",X"C2C4",X"CCC7",X"7DD1",X"FFE3",X"F6FA",X"F7F7",
      X"F8F8",X"FCF7",X"ABF1",X"FFDC",X"AEF6",X"FFC9",X"B3EB",X"FDE7",
      X"F4F3",X"F6F5",X"F6F5",X"F6F5",X"BFEE",X"B7ED",X"FDAD",X"F1F5",
      X"EEF1",X"EFEF",X"EBF9",X"DA9A",X"F3FE",X"EFEF",X"E7FA",X"D98C",
      X"F0FC",X"EEF0",X"E2F0",X"E6D1",X"A7E6",X"F8DD",X"F0F2",X"EDEF",
      X"EBEC",X"F7EC",X"97D2",X"F7E0",X"ADEF",X"F9CB",X"EBED",X"EDED",
      X"ECEB",X"E9E9",X"D3F0",X"EFBD",X"91BD",X"8E8C",X"9495",X"9092",
      X"8D8F",X"C899",X"D3CD",X"D3D7",X"C9CD",X"CDCB",X"D0C8",X"D8D7",
      X"DADE",X"CFD5",X"C5C7",X"D1C9",X"8ED1",X"FEF5",X"F5F5",X"F6F7",
      X"F4F5",X"FBF5",X"AAEB",X"FFE2",X"ABEA",X"FFEA",X"BACD",X"F7FB",
      X"F2F4",X"F4F4",X"F4F3",X"F7F4",X"C3DB",X"9FF6",X"FFBB",X"F0F3",
      X"EAEF",X"EFED",X"DFFB",X"E591",X"F0FB",X"EEF0",X"D8F0",X"E283",
      X"EFFD",X"EEEF",X"EFF0",X"CEDF",X"B9E8",X"F6BE",X"EEF0",X"EBEE",
      X"EBEC",X"EDEB",X"A1F0",X"F4B7",X"C0EF",X"F4B9",X"EAEC",X"EBEC",
      X"EAEB",X"EAEC",X"EEED",X"BAC4",X"BAF4",X"9092",X"9395",X"9293",
      X"8F90",X"9C8F",X"D2CE",X"D4D5",X"CBCE",X"CECD",X"D2CE",X"D8D8",
      X"DFE1",X"D5DB",X"C9CE",X"D6CE",X"A1CF",X"FBFF",X"F5F5",X"F6F5",
      X"F5F5",X"FDF5",X"A7E2",X"FFF0",X"BBD5",X"F6FB",X"D5B0",X"F2FE",
      X"EBF3",X"F3F0",X"F4F4",X"FAF3",X"C9CF",X"9BF7",X"FFC9",X"F1F1",
      X"E5EE",X"F0EC",X"CBFA",X"F290",X"F1F6",X"E6F5",X"D5D7",X"CF70",
      X"EFFD",X"EEEF",X"F1EF",X"D6EC",X"CDD3",X"E8A7",X"ECF3",X"EBEB",
      X"EBEB",X"EBEB",X"C5F7",X"E69F",X"C4F3",X"EFA6",X"EBEE",X"EBEC",
      X"EBEC",X"EBEA",X"EDEB",X"A5E2",X"F9AE",X"97B8",X"9794",X"9296",
      X"8D90",X"8D8C",X"DAA3",X"D8DA",X"D3D7",X"CDCF",X"D9D5",X"DADB",
      X"E0E2",X"D9DE",X"CED2",X"DAD3",X"AACC",X"FBFF",X"F5F4",X"F4F5",
      X"F5F4",X"FFF5",X"AEE0",X"FEF3",X"D1BB",X"D9FF",X"EFAC",X"F3F8",
      X"E6E7",X"F2F2",X"F3F3",X"F8F2",X"D4C1",X"93F4",X"FCD3",X"F3EE",
      X"E1E9",X"EFEF",X"BEFA",X"F59A",X"F1F3",X"DDF9",X"D5CD",X"A25C",
      X"F4F7",X"ECF1",X"F0EC",X"E4ED",X"C8CE",X"CE98",X"EFFA",X"EAEB",
      X"EAEB",X"EBE8",X"E9F0",X"CBA6",X"CEF6",X"E696",X"ECEF",X"EBEC",
      X"EAE8",X"EAE9",X"E9EE",X"CCCA",X"B38D",X"BDFB",X"96A0",X"9696",
      X"8E93",X"928E",X"A696",X"DEDC",X"D8DD",X"D0D3",X"DBD8",X"DDDD",
      X"E1E0",X"DBDF",X"D1D4",X"DDD5",X"B6CA",X"F9FF",X"F5F7",X"F4F4",
      X"F4F4",X"FEF4",X"AFDD",X"EBF5",X"E9B2",X"C7FE",X"FBC2",X"EDF4",
      X"EADA",X"F0F3",X"EFF0",X"F2F4",X"E1B6",X"84EB",X"FBDB",X"F5F0",
      X"DFE1",X"EEF0",X"AAFA",X"FCA7",X"F0F4",X"CDF9",X"CDCF",X"8E81",
      X"FBD3",X"EDF3",X"EEEA",X"EDEE",X"C3D8",X"A897",X"F1F8",X"EAEC",
      X"E9E9",X"E8EA",X"F7EB",X"A4BD",X"E2EF",X"D89C",X"ECF2",X"ECEC",
      X"E8E9",X"E7E8",X"EEEA",X"BFBC",X"71D3",X"FFBE",X"91B7",X"9696",
      X"9396",X"9694",X"9395",X"DEA0",X"D9DE",X"D4D5",X"DBD9",X"DBDA",
      X"E1DF",X"DCE0",X"D3D7",X"DFD8",X"BABB",X"F8FF",X"F4F6",X"F3F4",
      X"F4F4",X"FFF3",X"ADD8",X"D7F9",X"FAC1",X"B6F5",X"FCD6",X"E2F1",
      X"EED8",X"EFF0",X"EFEF",X"E6F6",X"EFAE",X"8BE4",X"F9E8",X"F2F1",
      X"DCD8",X"EFF2",X"9AF3",X"FCB6",X"EEEE",X"B0F3",X"B6C5",X"A999",
      X"EB96",X"EFFA",X"EDED",X"EEEB",X"D0E9",X"89A4",X"F5E8",X"EAEC",
      X"E8E8",X"E7EA",X"F0E8",X"9EDD",X"F0DD",X"C7A3",X"EBF4",X"EBEA",
      X"E7E7",X"E7E6",X"EEE8",X"9ED8",X"B9E3",X"D464",X"B0FE",X"948E",
      X"9495",X"9191",X"9495",X"A294",X"D4D9",X"D4D3",X"DAD9",X"D9D8",
      X"E1DF",X"D9DF",X"D2D4",X"DBD6",X"C4AD",X"F5FF",X"F3F5",X"F3F3",
      X"F3F3",X"FFF4",X"ABD5",X"C3F8",X"FDCC",X"ABE8",X"FBE4",X"D8EE",
      X"F1DE",X"EFF0",X"EFEF",X"D9F9",X"FDAD",X"8DCF",X"F7F4",X"EBF3",
      X"E3D2",X"F1F1",X"92E9",X"FACB",X"F0EA",X"9EEF",X"ACC8",X"DFB4",
      X"AB80",X"F3F9",X"EDED",X"EBED",X"EAEE",X"76BC",X"F9C9",X"ECEE",
      X"E7EB",X"E6E7",X"EBE7",X"B2EE",X"FACE",X"B4A8",X"EBF3",X"E7EA",
      X"E6DD",X"E6EA",X"EAE6",X"A6EE",X"EF8B",X"6394",X"FFD3",X"94BB",
      X"8A93",X"928B",X"9596",X"9696",X"CE9F",X"C5CB",X"DAD4",X"DFDF",
      X"DCDB",X"D6DB",X"CFD1",X"D3D0",X"C7A8",X"F4FF",X"F2F2",X"F3F3",
      X"F3F3",X"FEF3",X"B2D6",X"AFEC",X"FFE3",X"B5D2",X"F9F2",X"D1E3",
      X"F1E6",X"EFEF",X"EFEE",X"C7FA",X"FFB3",X"8DBF",X"F4F6",X"E3F2",
      X"E7CC",X"F4F0",X"8ADB",X"F6DB",X"F3EB",X"91DE",X"9CCD",X"F7C9",
      X"80BF",X"FBCB",X"ECF0",X"ECEC",X"F2ED",X"87DE",X"F5A9",X"EAEC",
      X"EAE9",X"E7E7",X"EAE9",X"C2EE",X"FAC2",X"ACAD",X"E9F1",X"E7EA",
      X"DECA",X"E5E8",X"E7E6",X"CBF2",X"A051",X"68EC",X"CF61",X"C6F9",
      X"8C98",X"908C",X"9290",X"9294",X"938E",X"C6B8",X"D2CF",X"D8D7",
      X"D8D9",X"D0D6",X"C9CB",X"CFCC",X"CDA6",X"F1FE",X"EFEF",X"F0F0",
      X"F3F3",X"FBF3",X"BAD8",X"AFD3",X"F7F5",X"C7B5",X"F2FB",X"D0D5",
      X"F0EC",X"EEEE",X"F2EE",X"B4F8",X"FFB6",X"94BA",X"F3F6",X"DAF2",
      X"EACC",X"F7EE",X"9CCF",X"F1EA",X"F9EC",X"8DCD",X"99CE",X"F8DD",
      X"AEEE",X"E292",X"ECF3",X"EAEA",X"ECEA",X"ABEE",X"EB8C",X"EBEE",
      X"E8E8",X"E8E5",X"E6E7",X"DBEB",X"EEB9",X"A4BD",X"E9EB",X"E8EA",
      X"D5BF",X"E4E7",X"E6E5",X"EBEB",X"7495",X"CDCE",X"A27B",X"E2BB",
      X"8DD0",X"8C97",X"928A",X"9295",X"8C8C",X"B38D",X"CECA",X"D4D3",
      X"D8DB",X"CED4",X"C9CA",X"CFCD",X"D1A7",X"F2FE",X"EDEE",X"EFEF",
      X"F2EF",X"FBF2",X"BADB",X"C0C0",X"EFF8",X"DBAB",X"E6F7",X"D4CA",
      X"EFF0",X"EDED",X"F2F2",X"A5E9",X"FFBE",X"9CB9",X"F1F8",X"D3F2",
      X"EACE",X"FAEE",X"9CBB",X"F0F1",X"F9EB",X"94B2",X"A6D3",X"F4EA",
      X"EAF5",X"A2A9",X"F3E4",X"E9EB",X"EAEB",X"D7F2",X"D17D",X"E9F0",
      X"E6E6",X"E7E6",X"E5E7",X"E8E7",X"DCC4",X"9BC4",X"EBE7",X"E7E7",
      X"D1BF",X"E1E6",X"E4E3",X"F0E6",X"9DC8",X"D1A1",X"ABB0",X"9E9D",
      X"D9D2",X"969D",X"928C",X"BEA7",X"8E95",X"8F8E",X"D2AF",X"D8D9",
      X"DCDB",X"D4D8",X"CED0",X"D3D0",X"D5B2",X"F2FD",X"EFEF",X"EFEF",
      X"EFEF",X"FCF1",X"A8D4",X"CCB0",X"E1FB",X"E6AC",X"DDF2",X"E1C6",
      X"EDF3",X"EEEE",X"CEF7",X"ABC0",X"FFD0",X"9FAB",X"F0F9",X"CBED",
      X"EAD0",X"F7EC",X"A3AD",X"EFF7",X"F8EB",X"9A90",X"B0C2",X"F4F5",
      X"F7F2",X"95E3",X"EB9F",X"E9F3",X"EBEB",X"EDEF",X"AD90",X"E9F1",
      X"E3E5",X"E6E6",X"E6E7",X"E9E7",X"D2D1",X"8AC5",X"EAE2",X"E9E5",
      X"C9B6",X"E0E8",X"E2E2",X"EDE3",X"A0D3",X"9EB2",X"99BF",X"9697",
      X"B09A",X"ADC7",X"9699",X"DDA4",X"A9D4",X"8E8E",X"B28F",X"DCDE",
      X"DCD9",X"DBDE",X"D4D7",X"D6D5",X"D9AF",X"F1FC",X"F1EF",X"F0EF",
      X"EEF0",X"FCEE",X"99D0",X"DBAE",X"D4FB",X"F0B6",X"D0EF",X"E9CA",
      X"EDF0",X"F3EC",X"9CF0",X"ADBA",X"FED5",X"AB9F",X"F0F8",X"C7E7",
      X"EBD1",X"EFEA",X"BCA6",X"EEF8",X"E4F1",X"AC70",X"BBAB",X"F3FA",
      X"F2F1",X"DBF6",X"A287",X"EDEB",X"E9EA",X"F2EC",X"96B5",X"EAED",
      X"E2E4",X"E5E3",X"E5E5",X"E7E5",X"D1DA",X"7BCC",X"EBDA",X"E7E5",
      X"BAB5",X"E4E9",X"E3E2",X"E9E3",X"A2E5",X"99A2",X"9FAB",X"989E",
      X"9494",X"B3A0",X"9FA1",X"C799",X"D9DC",X"9CBC",X"9493",X"D39F",
      X"DBD8",X"DDDF",X"D7D9",X"DAD8",X"DCB1",X"EFFC",X"EEED",X"EFED",
      X"ECEF",X"FAF0",X"92D5",X"EBB5",X"C1F9",X"F8BF",X"C7E6",X"EFD4",
      X"EDF0",X"F8EE",X"94DA",X"A2CA",X"FDDC",X"A087",X"EDF7",X"C3E2",
      X"E9D4",X"E6E8",X"C595",X"EEF8",X"BFF9",X"C258",X"D8A8",X"F2F9",
      X"EFF1",X"F8F1",X"87D3",X"F0B5",X"E9ED",X"F0EA",X"8ED4",X"EBDB",
      X"DFE4",X"E3E3",X"E5E3",X"E5E4",X"E0E1",X"8BD8",X"F1D4",X"EAE5",
      X"A7B3",X"E5E8",X"E4E2",X"E7E2",X"B9EC",X"949C",X"AFA2",X"97A5",
      X"9195",X"BC91",X"96AE",X"A7A0",X"DADD",X"D6D6",X"A1C6",X"9694",
      X"DCD9",X"DBDC",X"D5D7",X"DEDA",X"E6B1",X"EDFB",X"EDEB",X"EEEE",
      X"EDED",X"F6ED",X"92D9",X"F4CE",X"A2F0",X"F9CB",X"C3DD",X"EDDB",
      X"EDEE",X"F9EE",X"ADC5",X"91DE",X"F7E2",X"A364",X"E2F4",X"BBDA",
      X"E8D8",X"DCED",X"D38D",X"EEF5",X"8FFB",X"C657",X"EEA8",X"F1F7",
      X"EDF1",X"F3EE",X"CEF6",X"C38F",X"ECF4",X"EDE7",X"88E7",X"EAC2",
      X"E2E2",X"E4E4",X"E3E2",X"E2E2",X"E7E1",X"8FE2",X"EFC8",X"EBE5",
      X"90AA",X"E4DC",X"E5E0",X"D2E5",X"C7D4",X"979E",X"A09D",X"9B97",
      X"9595",X"A894",X"CDE4",X"92A5",X"9B81",X"D5CD",X"DCDB",X"A2C5",
      X"DCE0",X"D5D8",X"CDD0",X"D6D1",X"E8B5",X"ECFC",X"ECE9",X"EDED",
      X"EDED",X"F3ED",X"9DDE",X"F8DE",X"9FE0",X"F7E5",X"C2D0",X"F0E4",
      X"EEEF",X"F4ED",X"CAAE",X"77DB",X"EEE0",X"AD4B",X"CFE9",X"B7D2",
      X"EDDA",X"CEF3",X"E89A",X"F3EE",X"69E7",X"B583",X"F8B5",X"F1F5",
      X"EFF0",X"F0F0",X"F5F0",X"94C4",X"F2D3",X"ECE9",X"9DEE",X"E9A5",
      X"D7CF",X"E3E7",X"E4E4",X"DFE2",X"E5E0",X"88E5",X"EFBA",X"EFE4",
      X"7DA5",X"E7CF",X"E3E3",X"C3EA",X"D2A1",X"92A6",X"9C97",X"9B8D",
      X"8F93",X"918E",X"DCD8",X"9EBD",X"7C96",X"6160",X"D287",X"DEDD",
      X"DBDF",X"D2D6",X"C8CE",X"CDC9",X"E8B8",X"EBF9",X"EBE9",X"EDEC",
      X"ECEC",X"EFEB",X"A2E4",X"FBDB",X"A7CF",X"EBF1",X"C6C4",X"F1EC",
      X"ECEC",X"DEF1",X"E798",X"6AB6",X"DDE3",X"A83B",X"C0D7",X"B7CD",
      X"EDDA",X"B6F3",X"F0A6",X"F6ED",X"71BF",X"A1A7",X"FBCB",X"F2F3",
      X"F3F2",X"F6F4",X"F6F5",X"B3F6",X"DA93",X"ECEF",X"B3EE",X"E78B",
      X"C4B1",X"E2EC",X"E2E2",X"DEE1",X"E4E0",X"90E7",X"EDAC",X"EDE4",
      X"7AAD",X"E1BA",X"E0E0",X"D3E6",X"C27A",X"8FB8",X"9694",X"869B",
      X"8E98",X"8D8E",X"D8CD",X"9BDC",X"BA8F",X"87A3",X"7181",X"DAB3",
      X"D4D8",X"CFD1",X"C8CA",X"CCC8",X"EBC0",X"EDF4",X"ECEB",X"ECEB",
      X"ECEB",X"EEEC",X"A1E8",X"FED3",X"A6C5",X"DFEE",X"CFBD",X"EDEF",
      X"EDEC",X"B1F3",X"EBA5",X"7E88",X"CCE9",X"A432",X"B9C2",X"B5CC",
      X"ECD9",X"A7ED",X"F3B9",X"ECEF",X"8FA2",X"9DA8",X"F9E3",X"F7F5",
      X"F1F5",X"E6EB",X"DCE0",X"C7D7",X"7F88",X"BEB0",X"BDC4",X"E07D",
      X"AAB1",X"E0EC",X"E1DF",X"DEE0",X"E1DE",X"98E8",X"E998",X"EAE2",
      X"73AF",X"D2A9",X"E3E5",X"E7E3",X"9880",X"98CA",X"9292",X"819B",
      X"8D9A",X"8B8E",X"D4B0",X"C0D8",X"988E",X"CAC9",X"CFCD",X"D6D2",
      X"D2D5",X"CFD0",X"C9CD",X"CCCA",X"EDB9",X"EBF3",X"EDEB",X"EDED",
      X"EBEC",X"EBEB",X"A9E9",X"FECB",X"B2B9",X"D5F4",X"DBBB",X"EAED",
      X"F5EC",X"8CE5",X"BDCA",X"9282",X"BCDF",X"AF39",X"B7BA",X"B4CA",
      X"EADB",X"A0E4",X"F1D2",X"DCF1",X"A698",X"A99D",X"E3E7",X"C9D3",
      X"B1BE",X"A9AA",X"B1A9",X"C3BB",X"9FC5",X"AA77",X"D5D1",X"CD83",
      X"96C3",X"E4E4",X"DFDE",X"DDDF",X"DFDD",X"9DED",X"E791",X"EAE0",
      X"71AE",X"C7A5",X"E0E6",X"ECE0",X"72A3",X"A5C9",X"9290",X"9292",
      X"977E",X"8D8D",X"D89E",X"D7DC",X"8E9F",X"CABB",X"D4CC",X"DADA",
      X"DADC",X"D4D6",X"CACF",X"CBC8",X"EDB1",X"ECF2",X"ECEC",X"EDED",
      X"E9E8",X"EAE9",X"B4EE",X"F9BA",X"BFB5",X"CBF6",X"E0BD",X"E9E9",
      X"FBED",X"7BB0",X"97DD",X"96A6",X"BCCF",X"B456",X"B7AF",X"B5C5",
      X"F1E0",X"A6CE",X"EDE6",X"B8F2",X"9E9F",X"8776",X"BFB6",X"C8C4",
      X"D6D0",X"E5DD",X"F2ED",X"F3F3",X"F8F8",X"99C5",X"E5C6",X"B894",
      X"94D4",X"E5DE",X"DEDE",X"DADC",X"DBDB",X"A8E7",X"E494",X"E8DC",
      X"74B2",X"B89B",X"DFE0",X"EADD",X"60C7",X"A8B9",X"9591",X"9997",
      X"9A7C",X"8D8E",X"DD96",X"DEE2",X"8EC4",X"C8A2",X"DAD0",X"E0DF",
      X"DEE0",X"D8DC",X"CDD2",X"CECD",X"F2A8",X"EEF4",X"EDEE",X"ECED",
      X"E9E9",X"E8E9",X"BFEF",X"F0B0",X"C1AB",X"C3F1",X"E5C2",X"E9E7",
      X"EBF5",X"9967",X"93C6",X"ACCF",X"BFCC",X"AD6B",X"A299",X"B9C6",
      X"F0E3",X"B9B3",X"EFF0",X"83E2",X"6177",X"B462",X"EFE2",X"F4F4",
      X"F8F6",X"F6F7",X"F5F5",X"F3F6",X"F4F0",X"C9F7",X"BD98",X"A5A0",
      X"8CDD",X"E6D0",X"DFDF",X"DCDD",X"DADA",X"A9DF",X"E59B",X"E6DC",
      X"7ABA",X"A897",X"E0D8",X"E5DB",X"5CDC",X"AF9B",X"9699",X"989A",
      X"8794",X"9192",X"C996",X"DFE1",X"9ED9",X"C78E",X"DDD6",X"E4E3",
      X"DCDB",X"DBDC",X"D2D6",X"D8D4",X"F5AC",X"E8EC",X"EDED",X"EDED",
      X"EAE8",X"E6EA",X"D3EF",X"E5A8",X"CBAA",X"BBEC",X"EACB",X"EAE9",
      X"ABF6",X"C750",X"B59D",X"B6EF",X"BAC5",X"AA7A",X"8F91",X"BEC1",
      X"E6E3",X"D3B8",X"F0EC",X"7DB2",X"7989",X"F5AB",X"F3F8",X"F3F2",
      X"F3F3",X"F2F3",X"F4F2",X"F3F3",X"F0F1",X"F9F6",X"97CE",X"9385",
      X"88DF",X"E8C2",X"DFDF",X"DCDD",X"D4DA",X"ACD8",X"E69C",X"E7DE",
      X"74B9",X"A19A",X"E0CE",X"E1DA",X"71E5",X"B987",X"969A",X"9996",
      X"839A",X"939D",X"C096",X"E0DF",X"C8DC",X"B792",X"DFDA",X"E3E2",
      X"DBD9",X"DCDC",X"D5D6",X"D6D7",X"F9A9",X"CDC9",X"ECEF",X"ECEC",
      X"E9E7",X"E9E8",X"E3F0",X"CBA2",X"D4AA",X"BDE6",X"EED3",X"F2E9",
      X"5FE4",X"BD80",X"EC9F",X"BCF8",X"A9BB",X"BA91",X"7D93",X"BCBC",
      X"E7E0",X"E5DE",X"E3EB",X"C39D",X"83B1",X"F9CD",X"F0F1",X"F2F1",
      X"F3F2",X"F4F4",X"F7F5",X"FBFB",X"F5F7",X"F6F4",X"DBFB",X"768A",
      X"8FDD",X"ECB4",X"DDE0",X"DCDC",X"D2DC",X"A9D1",X"E79B",X"E5DE",
      X"6CA5",X"9C9D",X"DEC5",X"DCDA",X"8FE2",X"B378",X"96A3",X"9794",
      X"9399",X"949B",X"B29A",X"E2DE",X"D9DF",X"A5A1",X"E0DC",X"E0E0",
      X"DBDA",X"D6DB",X"CED2",X"C4D3",X"FDAB",X"C9B0",X"ECF4",X"EAEA",
      X"E5E6",X"E6E6",X"EEEB",X"ADAA",X"DDAE",X"BBDD",X"F0D9",X"F8F3",
      X"61B0",X"A8A3",X"FCD6",X"C8FB",X"99B5",X"B4AD",X"6F83",X"BAB8",
      X"EAE1",X"E5E8",X"CAE7",X"E9A8",X"7B91",X"F9E8",X"EFF2",X"F1F0",
      X"F5F3",X"FBFA",X"E9F3",X"D4DE",X"CBC9",X"F3DC",X"FFFE",X"88D9",
      X"A3D1",X"ECA0",X"DBE2",X"DCDC",X"D3DB",X"A3CE",X"E990",X"D9DB",
      X"6899",X"98A0",X"DBBC",X"DAD8",X"98DD",X"B47D",X"96AE",X"9596",
      X"9490",X"9276",X"A097",X"DFDD",X"D9DF",X"8DB0",X"DBD8",X"DBDC",
      X"DADA",X"D1D7",X"CACB",X"C5CF",X"FABE",X"D6A7",X"ECF6",X"EAEB",
      X"E7E7",X"E6E5",X"F3EA",X"93B7",X"E3B4",X"BFD9",X"EEDC",X"BFEC",
      X"5F74",X"685B",X"A39F",X"96AC",X"8182",X"A7BF",X"696A",X"BAB6",
      X"E7E0",X"E5E6",X"A3E4",X"ECC4",X"9465",X"F4F9",X"F0EF",X"F3F2",
      X"F1F7",X"C2DC",X"B7B5",X"A2AB",X"B6A5",X"CEC3",X"D5D6",X"90CB",
      X"ADC8",X"E992",X"DDE2",X"D9DC",X"D2DB",X"A7C9",X"EB90",X"C0D1",
      X"5C9C",X"969D",X"D7AF",X"DBD8",X"9ADE",X"AC87",X"93B0",X"9296",
      X"8D8E",X"9460",X"A095",X"DCDD",X"D2D9",X"8DBF",X"D9BE",X"DADB",
      X"D8D9",X"CCD3",X"C4C5",X"C6C8",X"F5C5",X"CC97",X"EBF8",X"E8EB",
      X"E6E9",X"E5E6",X"F5E7",X"78D0",X"D9A5",X"A6BF",X"ADAD",X"578C",
      X"444D",X"8C53",X"999C",X"90A0",X"7368",X"B7CF",X"5156",X"BCB3",
      X"E5DF",X"EDE4",X"81C3",X"D1E7",X"CA5B",X"F1FA",X"F2F1",X"F4F6",
      X"ABCC",X"99A3",X"8794",X"5370",X"3F43",X"2F33",X"2E37",X"3C31",
      X"B7B7",X"E085",X"DDE1",X"D9DB",X"C9DA",X"AFBE",X"EB9E",X"B1C7",
      X"539A",X"9B9B",X"D4A7",X"DAD9",X"A2E0",X"A196",X"92A7",X"9094",
      X"898C",X"8475",X"9D91",X"D9DB",X"CAD1",X"8EC7",X"D5AB",X"D8DB",
      X"D6D8",X"CAD2",X"C5C4",X"C6C7",X"F4CC",X"C28E",X"ECEC",X"E6E7",
      X"E6E6",X"E7E5",X"F1E9",X"68E2",X"A369",X"988B",X"C1B5",X"9199",
      X"8395",X"FECE",X"FFFF",X"E8FD",X"7B9A",X"C6DB",X"3741",X"C1A7",
      X"E4DE",X"ECE7",X"A693",X"AAFF",X"F485",X"F2F7",X"F7F3",X"AFE3",
      X"B0A4",X"4882",X"1427",X"1B15",X"191F",X"1B1B",X"4E23",X"5869",
      X"C8A1",X"DA88",X"DBE4",X"DADA",X"C7DC",X"ACBB",X"EB9A",X"A9BC",
      X"4BA8",X"9B94",X"CCA1",X"DBDA",X"A8DB",X"A9B1",X"92A0",X"9096",
      X"898B",X"9992",X"9A94",X"D9DC",X"C9D1",X"A4C9",X"D7A1",X"DADC",
      X"DADA",X"D2D8",X"CBCD",X"AECF",X"F5DA",X"C19C",X"E7C7",X"E5EA",
      X"E5E5",X"E6E5",X"EDEB",X"79EF",X"C755",X"C3BF",X"E0E6",X"B7AB",
      X"AF89",X"FEFC",X"FEFC",X"FCFF",X"66A6",X"E1E3",X"263D",X"BF92",
      X"E2D8",X"CCEF",X"E190",X"8EF3",X"FBBD",X"F0F3",X"E2F4",X"BFAC",
      X"58C1",X"310C",X"5865",X"272F",X"2126",X"272A",X"BF36",X"A7FC",
      X"CE8E",X"D38C",X"DAE2",X"DADB",X"C6DB",X"ACBB",X"E99D",X"A2AD",
      X"38AE",X"9E86",X"C89A",X"D9DA",X"B7D9",X"9C8D",X"949C",X"9196",
      X"8C8D",X"B097",X"9AC2",X"DBDF",X"D1D6",X"BACF",X"DBA1",X"DEDF",
      X"DFDD",X"DBDF",X"D4D6",X"AED8",X"E8E8",X"C494",X"E1AB",X"E5EC",
      X"E5E5",X"E5E4",X"E4E4",X"A4F4",X"DC5C",X"CBCF",X"B8ED",X"93BE",
      X"E47F",X"E5F4",X"C8D6",X"DAC6",X"5794",X"F7E6",X"3A65",X"C07E",
      X"E9DB",X"95DE",X"FEC2",X"A7D7",X"F5EA",X"F1F0",X"E2F1",X"B6DB",
      X"1A3B",X"9E63",X"779E",X"1E3F",X"131B",X"3F3A",X"F058",X"9EF1",
      X"C88C",X"CD81",X"D8E1",X"D8D7",X"C0DB",X"B2B8",X"E9A0",X"A9A9",
      X"2BAB",X"A174",X"C295",X"D8DA",X"BCDC",X"9592",X"9492",X"9294",
      X"9091",X"CE93",X"9ED3",X"DEE0",X"D8DC",X"D1D5",X"DFC4",X"E1E1",
      X"E0DD",X"DFE3",X"D5D7",X"99D8",X"D1FD",X"D377",X"DDA6",X"E6F0",
      X"E4E5",X"E3E2",X"E6E2",X"CEF1",X"C667",X"D5D5",X"ABC3",X"89C9",
      X"EDD6",X"C1D4",X"BABE",X"A3A8",X"456E",X"FDCE",X"6C88",X"AB6C",
      X"DADA",X"8F8A",X"F7F2",X"E3E1",X"F2F7",X"F0F0",X"F7F1",X"3BB7",
      X"B656",X"77E4",X"4A2C",X"3758",X"3A20",X"6474",X"CD78",X"ABB5",
      X"C88D",X"C47D",X"D7E2",X"D9D8",X"BADA",X"B0B3",X"ECA3",X"A099",
      X"31AB",X"9B61",X"B58F",X"D9D5",X"B4DF",X"8A91",X"948D",X"9293",
      X"9292",X"D493",X"9ACF",X"DFE2",X"DBDD",X"D5D7",X"E0DC",X"E2E2",
      X"DFDC",X"DDE1",X"D2D5",X"A3CA",X"B8FF",X"DE63",X"D1AF",X"E6F0",
      X"E5E5",X"E0E1",X"E1E2",X"EAE1",X"9D83",X"C7DB",X"D0A4",X"90A4",
      X"83B1",X"606A",X"826A",X"A098",X"5182",X"FFBE",X"8EAF",X"666E",
      X"7287",X"D977",X"F1F8",X"F3F1",X"F0F2",X"F1F0",X"CFF8",X"9A67",
      X"FFEF",X"9AFF",X"4C20",X"777A",X"B188",X"59A6",X"B377",X"CDE0",
      X"C883",X"C179",X"D6E3",X"DAD6",X"B5D7",X"ADB2",X"EEAC",X"9477",
      X"43A7",X"9356",X"AF92",X"DAD1",X"A1DF",X"9796",X"979B",X"9494",
      X"9193",X"CC93",X"A2D8",X"DFE2",X"DADC",X"D5D8",X"E1DB",X"E1E2",
      X"DCD9",X"D6DC",X"CDCF",X"B59F",X"87FF",X"E655",X"C0B2",X"E7EF",
      X"E2E4",X"E0E1",X"DDE3",X"EABF",X"74B2",X"94BF",X"9399",X"1E37",
      X"0C14",X"1812",X"1918",X"2724",X"4535",X"F49B",X"C3E3",X"9FC0",
      X"739A",X"F6B6",X"F0F1",X"F0F1",X"F1F0",X"F5F1",X"AEED",X"FABF",
      X"E3FB",X"C4DC",X"2450",X"6B4A",X"998E",X"938C",X"EFCF",X"D5F6",
      X"C38C",X"C282",X"D6E4",X"DAD7",X"ADD6",X"A7AF",X"E6B8",X"955C",
      X"509B",X"8B54",X"A894",X"D9D0",X"97DD",X"949C",X"94AA",X"9695",
      X"8E91",X"BF92",X"A8DA",X"DBDE",X"D0D6",X"CCCE",X"DDD3",X"DEE0",
      X"D9D8",X"D1D7",X"C8CA",X"C3A1",X"52F9",X"EE54",X"B3BB",X"E7F1",
      X"E0E1",X"E1E1",X"E4E2",X"BFA5",X"7BE7",X"4670",X"1A35",X"3A18",
      X"7967",X"2449",X"2828",X"1F2E",X"1C16",X"742F",X"EBC8",X"F8F8",
      X"C1F9",X"E996",X"EEF2",X"F1EF",X"F1F1",X"F3F1",X"E5ED",X"F7F8",
      X"B3EA",X"A599",X"8291",X"AA94",X"D4BE",X"F9E8",X"CEFF",X"D59D",
      X"BB9C",X"B97F",X"D6E4",X"DBD7",X"A6D1",X"A4AC",X"DAC5",X"9743",
      X"5F8B",X"8156",X"9F90",X"DAD0",X"9EDB",X"9291",X"94A0",X"9394",
      X"8D8E",X"C48F",X"C6D5",X"DADC",X"CDD3",X"C8C9",X"D9D0",X"DCDD",
      X"D6D6",X"CFD4",X"C9C9",X"E494",X"2DD6",X"E74A",X"ABCF",X"E7E9",
      X"DFE0",X"DFDF",X"EBDF",X"7DA5",X"9DF5",X"2023",X"905A",X"CAB2",
      X"85AD",X"2957",X"2021",X"422E",X"3240",X"8477",X"CB8D",X"F4F2",
      X"F0F6",X"C1A1",X"EFF7",X"F1EF",X"F0F1",X"F1F0",X"F5F4",X"F2F2",
      X"ECF1",X"EEEE",X"FAF6",X"FFFD",X"FBFE",X"F8F8",X"C1FA",X"E098",
      X"B8A0",X"B98B",X"D6E2",X"DAD8",X"A2CD",X"ABAC",X"CBD0",X"9232",
      X"6B78",X"7D59",X"9B8C",X"DBCE",X"A6D6",X"918F",X"9192",X"8D91",
      X"8D8C",X"CB8F",X"D8D4",X"D9DC",X"CCD3",X"C7C8",X"D6CE",X"DDDB",
      X"D6D8",X"CDD3",X"C9CB",X"FF93",X"13A5",X"E141",X"9FE0",X"E6DC",
      X"E0E0",X"DCDD",X"EDDE",X"44BD",X"E5BE",X"1248",X"DD71",X"FFFF",
      X"26B0",X"462F",X"0E2D",X"6423",X"515E",X"FFDF",X"E8EA",X"F3F3",
      X"F9F3",X"9DD0",X"F5EA",X"F1F1",X"F1F1",X"F0F0",X"F0F1",X"F0F0",
      X"F5F2",X"F8F6",X"F7F7",X"F8F6",X"F5F8",X"F2F2",X"F0F4",X"F1F1",
      X"B39A",X"C199",X"D6DE",X"D8D7",X"9DC5",X"B1B0",X"BDDB",X"8F26",
      X"7876",X"7757",X"9D8F",X"DCCF",X"A6CC",X"8E8D",X"9191",X"8D90",
      X"8E8C",X"CE98",X"DBD7",X"DCDF",X"CED5",X"C9CA",X"D8CF",X"E0DD",
      X"D9DB",X"CED5",X"BACA",X"FD9E",X"6870",X"D03B",X"8CEF",X"EAC6",
      X"DDE1",X"DADD",X"EADC",X"44D7",X"F86C",X"30AD",X"7B33",X"FFE9",
      X"6AFD",X"7136",X"2B5E",X"8C4D",X"5761",X"FFE5",X"F7FB",X"F2F3",
      X"F5F1",X"93EF",X"F8BE",X"F0F1",X"F0F0",X"EEF0",X"EFEF",X"F1F0",
      X"F2F3",X"F3F2",X"F3F3",X"F3F3",X"F4F4",X"F2F3",X"F3F1",X"F2F7",
      X"AB95",X"C39C",X"D5DE",X"D6D6",X"9DC1",X"B7B5",X"AAE5",X"8D1E",
      X"8380",X"6F5E",X"9B8E",X"DFCB",X"98BE",X"8B8A",X"9594",X"9093",
      X"8E8E",X"CDA6",X"DBD8",X"DCDD",X"D1D6",X"CFD0",X"DAD3",X"E2DF",
      X"DFDD",X"D7DC",X"90D3",X"D6BE",X"C745",X"BF46",X"95FA",X"EBAD",
      X"DCDF",X"DBDD",X"E2DB",X"76E8",X"BB3B",X"86EB",X"6082",X"DE76",
      X"DBFF",X"4E59",X"8476",X"93A4",X"684A",X"F7D6",X"F3F5",X"F1F2",
      X"F3F0",X"AFFB",X"F39A",X"EFF3",X"EEEF",X"EFEE",X"EFEF",X"F1F0",
      X"F1F2",X"F2F1",X"F2F2",X"F2F2",X"F3F3",X"F1F3",X"F2F1",X"F4F4",
      X"A89F",X"C896",X"D5DD",X"D5D7",X"97BC",X"C2B7",X"98E7",X"8124",
      X"7D6E",X"6665",X"958D",X"DEC4",X"A1B8",X"9290",X"9796",X"9496",
      X"9193",X"D4AD",X"D9D6",X"DADA",X"D7D8",X"D6D5",X"DCD7",X"E4E1",
      X"DFDC",X"DCE0",X"57D5",X"87E1",X"DE56",X"B747",X"A0FE",X"E696",
      X"DBDD",X"DCDE",X"D8D5",X"9AF2",X"8549",X"B9DF",X"D9A4",X"ADA9",
      X"CBCF",X"3086",X"704A",X"8477",X"DBA9",X"F5F3",X"F3F3",X"F0F2",
      X"F2F0",X"D2F9",X"E489",X"EFF6",X"EEED",X"EEEE",X"EFEF",X"F0F0",
      X"F1F1",X"F1F1",X"F1F1",X"F1F1",X"F2F2",X"F1F1",X"F2F2",X"F7F5",
      X"9BB1",X"D091",X"D6DB",X"D7D7",X"93B5",X"D4C3",X"84E3",X"7A43",
      X"6F7A",X"6251",X"8F90",X"DAC3",X"9CAF",X"9793",X"9695",X"9797",
      X"9396",X"DCC5",X"DCDC",X"DEDE",X"DADC",X"D7D7",X"DFD9",X"E1E2",
      X"E0DB",X"DBE2",X"63A9",X"3ED3",X"E2B2",X"A257",X"9DFF",X"DE69",
      X"DCE1",X"DEDE",X"CFD2",X"B2EF",X"8861",X"DAA9",X"BF86",X"EFFE",
      X"D8E3",X"B7C5",X"CABD",X"ECD4",X"FCFC",X"F4F5",X"F2F1",X"F1F1",
      X"F0F0",X"ECF5",X"C88E",X"F1F9",X"EFF0",X"EFEE",X"F0EF",X"F1F0",
      X"F1F1",X"F0F1",X"F1F0",X"F1F1",X"F1F2",X"F2F1",X"F2F2",X"F9F4",
      X"8CB2",X"D598",X"D6DB",X"D7D7",X"96AA",X"DDCE",X"7DD4",X"6F5A",
      X"9DA5",X"5965",X"908D",X"CFC1",X"B3A0",X"98C1",X"9898",X"9998",
      X"9496",X"DCD3",X"E3E2",X"E3E4",X"DCE1",X"D4D8",X"E2DD",X"DFE1",
      X"DBDD",X"D8D9",X"8360",X"3F93",X"DFD9",X"8E63",X"A8FF",X"B943",
      X"DEE6",X"DCDD",X"C5D3",X"CAE2",X"AB65",X"C497",X"87B6",X"F9E8",
      X"F9F8",X"FDFC",X"FDFE",X"F6FA",X"F2F3",X"F1F1",X"F0F1",X"F0F1",
      X"EFEF",X"F7F2",X"B6AA",X"F1F7",X"F0F0",X"EFEF",X"EFEF",X"F1EF",
      X"F1F1",X"F0F0",X"F0F0",X"F1F1",X"F2F1",X"F2F2",X"F2F1",X"FBF4",
      X"81B2",X"DA96",X"D5DB",X"D1D5",X"9C9F",X"DFD3",X"7DBF",X"6D5E",
      X"9699",X"6C98",X"918C",X"B9C2",X"D09F",X"C1D1",X"9897",X"9899",
      X"9E95",X"D4CD",X"E1D9",X"E0E3",X"D4DC",X"D0CF",X"DEDA",X"DFE1",
      X"D8DA",X"C4D7",X"A942",X"7D4E",X"D9D8",X"7497",X"C3FD",X"9352",
      X"E1E3",X"DBDD",X"C3D5",X"DFCF",X"906B",X"92C9",X"95D1",X"F7AB",
      X"F4F5",X"F5F5",X"F4F5",X"F1F3",X"F0F0",X"EFF0",X"F0F0",X"EFF0",
      X"EEEF",X"F5F0",X"C4CE",X"F1F3",X"F0EF",X"F0F0",X"EFEF",X"F0F0",
      X"F1F1",X"F0F0",X"F1F0",X"EFF0",X"F1F0",X"F1F1",X"F2F2",X"FDF4",
      X"6BBA",X"E08B",X"D4DB",X"C9D3",X"A596",X"E1D7",X"8BA7",X"6F5E",
      X"9295",X"8193",X"9A8F",X"93A1",X"CDA0",X"CBCD",X"9595",X"9394",
      X"BA92",X"CBC9",X"DBD4",X"DBDD",X"CDD5",X"CECC",X"D8D3",X"DDDD",
      X"D5D7",X"A3D4",X"9957",X"C638",X"D5D1",X"67B4",X"CEF8",X"8F8E",
      X"E4D2",X"DADB",X"C5D9",X"E8BD",X"5098",X"A9D0",X"C39D",X"CB81",
      X"F5FA",X"F4F3",X"F0F3",X"EFEF",X"EFEF",X"EFF0",X"EFEF",X"EFEE",
      X"EFEF",X"F0EF",X"E5E7",X"EEF1",X"F0EF",X"F1F1",X"F0EF",X"F0F1",
      X"F0F0",X"F0F1",X"F1F1",X"EEF0",X"F0EF",X"F2F1",X"F2F2",X"FAF4",
      X"5EBE",X"E586",X"D2D9",X"BFD5",X"B08D",X"DADA",X"B393",X"816A",
      X"9193",X"8491",X"7C7B",X"968F",X"CCA8",X"C6CA",X"9291",X"998F",
      X"C9BE",X"C6C6",X"D6CF",X"D5D8",X"C9D2",X"CCC8",X"D4CE",X"DBDA",
      X"D5D8",X"6CD4",X"5D7F",X"C980",X"D4CF",X"5DB8",X"CCEA",X"97A4",
      X"E8B6",X"DADD",X"CAD7",X"D6B3",X"42C3",X"E080",X"AF8F",X"8AAB",
      X"FAE2",X"F3F5",X"F0F1",X"EEEF",X"EFEE",X"EFF0",X"EEEE",X"EFEE",
      X"EFEF",X"F0EF",X"F5F3",X"EEF3",X"F0EE",X"EFF0",X"F0F0",X"F1F1",
      X"F0F0",X"F0F0",X"EFEF",X"EEF0",X"F0EE",X"F1F1",X"F2F2",X"FAF4",
      X"4EB8",X"E482",X"D1D7",X"B7D9",X"BA89",X"CDDE",X"A186",X"9B77",
      X"9295",X"8490",X"9974",X"93B7",X"CBBB",X"C7C9",X"928F",X"CBB2",
      X"C9CB",X"C9C9",X"D8D1",X"D9DB",X"CDD4",X"CECA",X"D6D0",X"DCDC",
      X"D8DC",X"57D3",X"4780",X"CEC8",X"DAD2",X"4FD5",X"CFD2",X"B8A0",
      X"DF9A",X"DADF",X"D2D6",X"BDB3",X"76DD",X"C059",X"82DB",X"9DB7",
      X"F498",X"F3F8",X"F1F0",X"EFEF",X"EFED",X"EFF0",X"EFEF",X"EFEE",
      X"EFEF",X"EFEF",X"EDF1",X"F2EC",X"F1EF",X"EFEE",X"F0F0",X"F1F1",
      X"F0F0",X"F1F1",X"EFEF",X"EFF0",X"F0EF",X"F1F1",X"F2F2",X"FCF6",
      X"31A1",X"E27F",X"D5D7",X"A6D6",X"C491",X"B4DE",X"9082",X"9590",
      X"9696",X"9594",X"9F96",X"A1D4",X"CFCF",X"CECE",X"CFAF",X"D1D9",
      X"CBCC",X"CFCA",X"DED6",X"DEDF",X"D2DA",X"D1CE",X"DAD5",X"E0E0",
      X"DCE0",X"639E",X"8E56",X"D5D2",X"E1DB",X"40E0",X"DAB3",X"D29C",
      X"CC9C",X"D9E0",X"D6D6",X"A8BF",X"A4DC",X"906B",X"C7EA",X"BA82",
      X"B593",X"F5F8",X"F1F2",X"F0F1",X"EFEF",X"EFF0",X"EFF0",X"EFEE",
      X"EFF0",X"EFEF",X"D0F5",X"F5BC",X"F1F4",X"F0EF",X"F1F2",X"F1F1",
      X"F0F1",X"F1F1",X"F1F0",X"EFF2",X"F0EF",X"F0EF",X"F3F1",X"FBF7",
      X"2B89",X"DD78",X"D5DA",X"9ACE",X"CA9A",X"9ADA",X"9488",X"969C",
      X"9698",X"9596",X"AD97",X"B2D5",X"D1D4",X"D5D2",X"E1DB",X"D9E0",
      X"CDD3",X"D4CE",X"DFD9",X"DFE0",X"D7DE",X"D4D2",X"DCD8",X"E3E1",
      X"DEE2",X"5C4A",X"CF4B",X"DAD6",X"E2E0",X"6ED9",X"E086",X"D88D",
      X"B2C7",X"DAE0",X"D6D7",X"A4CD",X"C9C4",X"8D7A",X"FAAF",X"8AAC",
      X"8FB9",X"F6C3",X"F1F3",X"F1F1",X"F0F0",X"F0F0",X"EFEF",X"EFEE",
      X"F0F0",X"EEEE",X"D8F7",X"E393",X"F0F8",X"F0F0",X"F0F0",X"F1F1",
      X"F1F1",X"F0F0",X"F0F1",X"EEF0",X"F0EF",X"F0F0",X"F2F1",X"F5F8",
      X"5B7B",X"D27C",X"D4DC",X"91C5",X"CCA4",X"89D7",X"928B",X"9598",
      X"9695",X"9596",X"BF99",X"D4DD",X"D4D7",X"DAD6",X"E2E0",X"DCE0",
      X"D2D8",X"D8D3",X"DFDB",X"DEDE",X"DBDF",X"D7D6",X"DEDA",X"E4E1",
      X"CBE1",X"4241",X"D7B3",X"DCD8",X"DFE0",X"7FC2",X"DD65",X"D992",
      X"A5DD",X"DCD5",X"D7D9",X"B0D6",X"D6A9",X"928D",X"CE99",X"B0FB",
      X"AA95",X"D395",X"F3F9",X"F0F1",X"EFF0",X"F0EF",X"EFEF",X"F0EF",
      X"EFF0",X"EEEE",X"F1F3",X"C79F",X"F0FA",X"F0F0",X"EEED",X"F0EF",
      X"F0F0",X"F0EF",X"EFEF",X"EFF0",X"F1EF",X"F1F1",X"F3F1",X"ECFB",
      X"967F",X"C983",X"D1DC",X"8CB6",X"D8B2",X"7CBE",X"9492",X"9395",
      X"9292",X"9493",X"DA98",X"DEDF",X"D7D8",X"DCD8",X"DFE0",X"DBDD",
      X"D7DD",X"DBD7",X"DFDF",X"DDDD",X"DDDF",X"DCDB",X"DFDC",X"E4E1",
      X"94E4",X"9A33",X"CCD0",X"D6D1",X"DCDB",X"9BAC",X"CD49",X"CCA6",
      X"C0DB",X"DFB9",X"D5D9",X"C1D6",X"C69E",X"90AF",X"9DBC",X"FCF3",
      X"96BA",X"9797",X"FAE0",X"F1F4",X"EFF0",X"F0EF",X"F0EF",X"F0F0",
      X"F0EF",X"EFF0",X"F5F1",X"BCC2",X"F1F7",X"F0EF",X"F0F0",X"EFEF",
      X"F0EF",X"F0F0",X"EFF0",X"F0F0",X"F0F0",X"F1F1",X"F3F2",X"DEFB",
      X"C299",X"CB88",X"CED8",X"94A9",X"C0B7",X"9097",X"918C",X"9393",
      X"9795",X"9194",X"E3C1",X"D7DF",X"CCD0",X"D6D1",X"DCDB",X"E0DF",
      X"D3DA",X"D3D1",X"DEDB",X"DFE0",X"D7DC",X"D4D5",X"DFDB",X"DDE0",
      X"36DD",X"D341",X"CBCB",X"D3CE",X"D7D8",X"8F96",X"B33A",X"C1AE",
      X"D7D4",X"D5A6",X"D5DC",X"CDD4",X"A0A7",X"8BC2",X"A8CA",X"FEBC",
      X"D0FA",X"80A0",X"E899",X"F5FC",X"EEF0",X"F0F0",X"EFEF",X"F0F0",
      X"F0F0",X"F0F0",X"F1F0",X"D7E4",X"F2F3",X"F0EF",X"F1F1",X"F0F1",
      X"F0F0",X"F1F0",X"EFF0",X"F0F0",X"F0F0",X"F2F1",X"F5F3",X"D7F9",
      X"D1C5",X"CA86",X"CBD7",X"8C9D",X"9BB1",X"8D91",X"8E8C",X"9290",
      X"9F93",X"CAB8",X"DDDE",X"D4DA",X"CBCB",X"D3CE",X"DAD8",X"DADC",
      X"CDD5",X"CECD",X"D9D4",X"D9DC",X"CED3",X"CDCC",X"D5D3",X"DCDA",
      X"57B6",X"CEC3",X"C7C9",X"D2CD",X"B1D5",X"C799",X"8B58",X"ACBB",
      X"D2CB",X"B3B7",X"D9DF",X"D3D4",X"78BB",X"A3A4",X"D696",X"E1A0",
      X"FDFC",X"9EDF",X"886E",X"FBE0",X"F0F5",X"EFF0",X"EFEF",X"F1EF",
      X"F1F1",X"F1F0",X"F1EF",X"EFF1",X"F1F0",X"F0F1",X"F1F1",X"F0F0",
      X"F0F0",X"F0EF",X"EFF0",X"F0F0",X"F1F1",X"F2F2",X"F4F3",X"DDF4",
      X"C8EA",X"CB75",X"ABD7",X"956F",X"8E92",X"8D8D",X"8C8C",X"918D",
      X"D6A2",X"CCD2",X"D8D7",X"CED4",X"C7C9",X"D2CD",X"D9D5",X"D4D8",
      X"C9CE",X"C8C7",X"D2CB",X"D5D8",X"C9CE",X"CECA",X"CDCB",X"DDD6",
      X"D5D4",X"CED4",X"C8CA",X"D0CD",X"D4D3",X"D1D8",X"57A4",X"A0BE",
      X"D4CD",X"90D3",X"DDD3",X"D1D6",X"89CB",X"B15F",X"9A6C",X"B5A6",
      X"FBF9",X"E6F9",X"5CAD",X"CA67",X"F7F5",X"F1F2",X"EEEE",X"F0EF",
      X"F0F0",X"EFF0",X"F2F0",X"EFF1",X"F0EF",X"F0F1",X"F0F0",X"EFF0",
      X"EFF0",X"EFEF",X"EFF0",X"F1F0",X"F0F1",X"F3F1",X"F3F3",X"EDF2",
      X"B6FD",X"C068",X"80A4",X"988A",X"8F92",X"8D8B",X"8C8D",X"A38D",
      X"D8D3",X"CBD2",X"D5D5",X"CED4",X"C8CA",X"D0CD",X"D9D3",X"D1D8",
      X"CACD",X"C9C8",X"D4CD",X"D8D8",X"CED3",X"CECD",X"D0CD",X"DED9",
      X"D9D9",X"D2D7",X"CDCD",X"D4D0",X"DCD5",X"D4DB",X"42C6",X"96AA",
      X"DCD2",X"B3DF",X"DFB4",X"D1D6",X"B4D2",X"875B",X"3690",X"6867",
      X"FDC3",X"F7F7",X"D7F9",X"909F",X"DDB0",X"F0EF",X"EEEE",X"EFEF",
      X"EFEF",X"EFEF",X"F0EF",X"F0F0",X"F0EF",X"F0F0",X"EFEF",X"EFEE",
      X"EEEF",X"F0EE",X"F0F1",X"F1F0",X"EFF0",X"F2F2",X"F3F3",X"F7F2",
      X"9BFE",X"8145",X"9995",X"9693",X"9293",X"8D91",X"A18D",X"D7CA",
      X"DCDD",X"D3D7",X"D9D9",X"D2D7",X"CDCD",X"D4D0",X"DCD5",X"D4DB",
      X"D0D1",X"CECD",X"DCD9",X"DEDF",X"D5DA",X"CDD0",X"D9D4",X"DFDE",
      X"DDDD",X"D8DB",X"D3D4",X"D6D5",X"E0D9",X"D9DF",X"62D8",X"9A7F",
      X"DEC8",X"DDDF",X"CBA1",X"CFD8",X"C7D0",X"5488",X"5CA4",X"364A",
      X"DC58",X"F3FD",X"F7F4",X"E5F8",X"BEC8",X"EDDA",X"EEED",X"EEEE",
      X"EFEF",X"EEEE",X"EEEE",X"EFEE",X"EFF0",X"EFF0",X"EFF0",X"EFEE",
      X"EEEE",X"EEEC",X"F0EF",X"F0F0",X"F0F0",X"F2F2",X"F3F1",X"FEF4",
      X"51EA",X"983B",X"968F",X"9498",X"9693",X"9095",X"DAB4",X"DBDE",
      X"DEDD",X"DBDC",X"DDDD",X"D8DB",X"D3D4",X"D6D5",X"E0D9",X"D9DF",
      X"D5D8",X"D8D3",X"DEDE",X"E0DF",X"DBDF",X"D0D4",X"DFD9",X"E0E0",
      X"DFDE",X"D9DF",X"D7D8",X"DAD8",X"E4DE",X"DEE1",X"A6DF",X"A24E",
      X"DEAC",X"DFDE",X"ADC9",X"D4DA",X"CECF",X"5CB5",X"8E5F",X"7C69",
      X"7E52",X"F8F0",X"F0F0",X"F5F2",X"EFF6",X"EFEC",X"EEED",X"EEEE",
      X"EFEE",X"EEEE",X"EEEE",X"EEEE",X"EFEF",X"F0F0",X"F0F0",X"EEF0",
      X"EDED",X"EEED",X"F0F0",X"F0F0",X"F1F0",X"F2F2",X"F4F2",X"FEF9",
      X"1C97",X"918D",X"9892",X"9497",X"9894",X"A598",X"DDD6",X"DEE1",
      X"DEDD",X"DCDC",X"DFDE",X"D9DF",X"D7D8",X"DAD8",X"E4DE",X"DEE1",
      X"D8DF",X"DCD5",X"DEDE",X"DFDE",X"DEE0",X"D6D8",X"E1DD",X"E2E1",
      X"DFDE",X"DBDE",X"D9D9",X"DDDA",X"E5E0",X"E1E3",X"CEE1",X"8C35",
      X"E093",X"E0E0",X"A9DF",X"D9BF",X"D1D4",X"87CB",X"6C2E",X"8170",
      X"5094",X"FA9E",X"EFF3",X"F1EF",X"F1F1",X"F0F1",X"ECEE",X"EEED",
      X"EEEE",X"EEEE",X"F0EF",X"EEEE",X"EEEE",X"EFEF",X"F0F0",X"EEF0",
      X"EEEC",X"EFEF",X"F0EF",X"F0F1",X"F2F1",X"F2F2",X"F7F2",X"CAFE",
      X"2641",X"91A1",X"9594",X"9596",X"9793",X"AF99",X"DCD9",X"E2E0",
      X"DCDD",X"D9DA",X"DFDE",X"DBDE",X"D9D9",X"DDDA",X"E5E0",X"E1E3",
      X"D9E1",X"DED5",X"E1E1",X"E0E0",X"DCDF",X"D7D8",X"E0DE",X"E2E1",
      X"DCDE",X"D8DC",X"D4D5",X"D8D6",X"E0DF",X"DEE4",X"D4D3",X"6261",
      X"CF90",X"E1E2",X"CBDA",X"D0A2",X"D4D5",X"B4D4",X"2E4B",X"5C5F",
      X"7F94",X"C64F",X"F1FA",X"EFEF",X"EFEF",X"EFEE",X"EDEF",X"EDEE",
      X"EEEE",X"EFEF",X"F1F0",X"EEF1",X"EEEF",X"EFEE",X"F0EF",X"EFF0",
      X"F1F1",X"EFEE",X"F0EE",X"F1F1",X"F2F1",X"F3F3",X"FCF4",X"85D6",
      X"224A",X"9653",X"9296",X"9794",X"9498",X"9292",X"CFA8",X"DED8",
      X"DBE0",X"D1D6",X"DCDE",X"D8DC",X"D4D5",X"D8D6",X"E0DF",X"DEE4",
      X"D4D3",X"D7D8",X"DEDB",X"E1E2",X"D9DA",X"D2D8",X"DDD5",X"E1E3",
      X"DCDB",X"D6DA",X"D0D1",X"D4D2",X"DAD9",X"D8DC",X"D0D1",X"49C0",
      X"B17E",X"DFE1",X"D2D7",X"B1C0",X"D4D5",X"CECF",X"327B",X"4E4B",
      X"9764",X"6B65",X"F8E2",X"F0F0",X"EDEF",X"EEEE",X"EEEF",X"EDEE",
      X"EFEE",X"F1F1",X"F5F4",X"F4F5",X"F1F2",X"EEF0",X"EEF0",X"E8EC",
      X"C2DC",X"ECC9",X"F0F1",X"F0F0",X"F2F1",X"F6F4",X"DCFB",X"A589",
      X"1D66",X"2420",X"8F7D",X"9591",X"9095",X"8E8D",X"968E",X"D9D2",
      X"D8DF",X"CBD1",X"DCDB",X"D6DA",X"D0D1",X"D4D2",X"DAD9",X"D8DC",
      X"D0D1",X"D5D5",X"DEDC",X"DFE1",X"D2D7",X"CBD0",X"D7CE",X"DADC",
      X"DAD9",X"D4D8",X"CBCD",X"D0CC",X"D5D3",X"D4D6",X"CDCC",X"8FD1",
      X"8564",X"DADA",X"CED3",X"9FCF",X"D5B6",X"D3CE",X"4FB2",X"4F52",
      X"714A",X"4071",X"EC8F",X"F1F8",X"EEF0",X"EDEC",X"EEEE",X"EDEE",
      X"EEED",X"F0EF",X"B4D0",X"CCBE",X"E8DA",X"EFEF",X"E0EB",X"C8D3",
      X"C7C2",X"F2E0",X"F0F0",X"EFEF",X"F2F1",X"FDF6",X"98DC",X"D3AE",
      X"1C60",X"1B28",X"9634",X"948E",X"9194",X"8D8E",X"8D8D",X"D8BD",
      X"D5DA",X"C9CE",X"DAD9",X"D4D8",X"CBCD",X"D0CC",X"D5D3",X"D4D6",
      X"CDCC",X"D2D1",X"D8D4",X"DADC",X"CED3",X"CBCF",X"D2CD",X"D9D7",
      X"DAD9",X"D2D8",X"C8CA",X"CFCA",X"D5D2",X"D4D6",X"CECF",X"CDCE",
      X"6376",X"D8BF",X"D0D4",X"C9CF",X"CB8E",X"D3D6",X"79D7",X"695A",
      X"4449",X"975A",X"9C93",X"FAEB",X"EEF3",X"EDED",X"EFEE",X"EEEF",
      X"EEEE",X"EEEE",X"C0DA",X"C1B5",X"E3D4",X"EFED",X"E9ED",X"E8E4",
      X"F2EC",X"F1F5",X"F0F0",X"F0F0",X"F5F3",X"D6FC",X"AD8F",X"D2D9",
      X"1D5D",X"2228",X"9220",X"948E",X"9294",X"9191",X"9090",X"DAAC",
      X"D4D8",X"CDD0",X"DAD9",X"D2D8",X"C8CA",X"CFCA",X"D5D2",X"D4D6",
      X"CECF",X"D2CE",X"D5D0",X"D8DA",X"D0D4",X"D0CF",X"D3D0",X"DAD7",
      X"DDDC",X"D4D9",X"C9CC",X"D3CF",X"DBD8",X"D9DC",X"D0D5",X"D0CF",
      X"7ECF",X"DB69",X"D0D6",X"D1CF",X"A0B6",X"D7D8",X"B4DB",X"7457",
      X"1F53",X"B164",X"8C9C",X"E68F",X"F2FA",X"EEEF",X"EFEF",X"EFF0",
      X"EEEF",X"EFEE",X"F5F1",X"F2F4",X"ECEF",X"EEED",X"F0EE",X"F2F1",
      X"EDF0",X"EFED",X"F0EF",X"F3F3",X"FBF6",X"8FDA",X"D1A9",X"CED7",
      X"215B",X"2729",X"821C",X"9591",X"9393",X"8F91",X"918F",X"DC9F",
      X"D8DB",X"D3D6",X"DDDC",X"D4D9",X"C9CC",X"D3CF",X"DBD8",X"D9DC",
      X"D0D5",X"D0CF",X"DCD8",X"DCDF",X"D0D6",X"D1CF",X"D5D4",X"DBD8",
      X"DFDF",X"D6DC",X"D0D1",X"D8D4",X"E0DD",X"DEE0",X"D4DB",X"D4D2",
      X"DEDF",X"8F62",X"D5DC",X"D4D2",X"A3DC",X"D8B2",X"D7D4",X"4980",
      X"7067",X"9A3D",X"9698",X"9198",X"F7CF",X"F0F4",X"EFEF",X"EEEE",
      X"EFEE",X"EEEE",X"F0EE",X"EEEF",X"EFEF",X"EFEF",X"EDED",X"EEEE",
      X"EDEE",X"EEEE",X"EFEF",X"F5F2",X"D4FB",X"AD98",X"CFD1",X"C9D5",
      X"2054",X"2A24",X"5D21",X"9697",X"9695",X"8F94",X"918E",X"DD98",
      X"DEE0",X"D8DA",X"DFDF",X"D6DC",X"D0D1",X"D8D4",X"E0DD",X"DEE0",
      X"D4DB",X"D4D2",X"E3DF",X"E1E4",X"D5DC",X"D4D2",X"DCDC",X"DFDF",
      X"E0DF",X"DCDF",X"D6D8",X"DCD8",X"E0DF",X"DFDF",X"D8DC",X"D9D6",
      X"E3DF",X"80DC",X"DAC0",X"DBD8",X"DDE0",X"BC90",X"D9D7",X"4EC0",
      X"DEA5",X"4CB5",X"989F",X"9A97",X"B882",X"F6F3",X"EEEF",X"EFEE",
      X"EEEE",X"EFEF",X"EEEE",X"EDED",X"EEEE",X"EDEE",X"EEEE",X"EEEE",
      X"EEEF",X"EFEF",X"F1EF",X"FBF5",X"87CA",X"D3AB",X"CBCF",X"CBD2",
      X"1C59",X"2A1F",X"2E29",X"96A2",X"9795",X"9196",X"9391",X"C196",
      X"DFE0",X"DCDC",X"E0DF",X"DCDF",X"D6D8",X"DCD8",X"E0DF",X"DFDF",
      X"D8DC",X"D9D6",X"E3DF",X"E2E2",X"DAE1",X"DBD8",X"E2E0",X"E1E1",
      X"E0DF",X"DDE0",X"DBDC",X"DEDD",X"E0DE",X"DBDC",X"D8DC",X"DED7",
      X"E4E0",X"E4E3",X"D8CE",X"DDD9",X"E0DE",X"81CB",X"D7B9",X"8ADB",
      X"E0A0",X"B1E5",X"9B83",X"9698",X"8998",X"DC9A",X"F6F7",X"EEF1",
      X"EEEE",X"F0EF",X"EFF0",X"EEEE",X"EEEF",X"EEEE",X"EFEF",X"EEEF",
      X"EFF0",X"EFEF",X"F6F1",X"C2F9",X"A67C",X"CFD1",X"CBCB",X"CFD1",
      X"1A63",X"2C20",X"172E",X"966F",X"9891",X"9597",X"9593",X"9B96",
      X"DCDC",X"DFDE",X"E0DF",X"DDE0",X"DBDC",X"DEDD",X"E0DE",X"DBDC",
      X"D8DC",X"DED7",X"E4E0",X"E4E3",X"DCE3",X"DDD9",X"E0DE",X"DEDE",
      X"DFE1",X"DADE",X"D3D6",X"DBD6",X"DFD9",X"DADF",X"D0D4",X"D5D0",
      X"E0DE",X"E4E4",X"D8DE",X"D1D4",X"DBD8",X"BFDE",X"9768",X"B8CC",
      X"D57A",X"E0DC",X"98BA",X"9493",X"9292",X"8AB1",X"EEBB",X"F2F6",
      X"EEEF",X"F0EF",X"F0F1",X"EFF0",X"EFEF",X"EFEF",X"F1F0",X"F0F1",
      X"EFF0",X"F0EF",X"F7F7",X"7EB6",X"CFAA",X"CACD",X"CCCC",X"D3D2",
      X"1F6E",X"2B26",X"202D",X"9A20",X"9296",X"9290",X"9193",X"9390",
      X"DCB4",X"DFDE",X"DFE1",X"DADE",X"D3D6",X"DBD6",X"DFD9",X"DADF",
      X"D0D4",X"D5D0",X"E0DE",X"E4E4",X"D8DE",X"D1D4",X"DBD8",X"E0DE",
      X"DDDF",X"D7D9",X"CDD1",X"D5D0",X"DBD6",X"D8DB",X"CDD3",X"D1CC",
      X"DBD9",X"DDDE",X"D4D8",X"D0D1",X"D6D3",X"DFDC",X"9DCA",X"B2A9",
      X"8B76",X"DFD9",X"C0DF",X"9AA0",X"8E8E",X"D299",X"8D9D",X"F3C7",
      X"F3F6",X"F1F1",X"F1F1",X"F1F1",X"F1F1",X"EFF0",X"F1EF",X"F1F1",
      X"EFF0",X"F7F1",X"ACF0",X"B483",X"CACF",X"CAC9",X"CCCC",X"D5D6",
      X"2774",X"2B2A",X"292B",X"4E16",X"909B",X"8E8E",X"8E8F",X"938F",
      X"D297",X"CDD3",X"DDDF",X"D7D9",X"CDD1",X"D5D0",X"DBD6",X"D8DB",
      X"CDD3",X"D1CC",X"DBD9",X"DDDE",X"D4D8",X"D0D1",X"D6D3",X"DFDC",
      X"D7DA",X"D2D6",X"C7CC",X"CFCA",X"D8D1",X"D5D9",X"CDD0",X"CDC9",
      X"D6D4",X"D8D8",X"D0D4",X"CDCD",X"D2CD",X"DFDB",X"D0DA",X"CBCB",
      X"A5B8",X"DCD5",X"D4DB",X"CCCE",X"A7B8",X"D19F",X"BDDD",X"AA91",
      X"F8D8",X"F6FC",X"F1F2",X"F2F2",X"F1F2",X"F1F0",X"F1F1",X"F3F1",
      X"F2F1",X"E8F8",X"91A7",X"CEBB",X"C8C9",X"CAC9",X"D1CC",X"B5E0",
      X"2B3F",X"292E",X"2A2B",X"1623",X"9084",X"8C8C",X"8D8C",X"918E",
      X"A396",X"CAD0",X"D7DA",X"D2D6",X"C7CC",X"CFCA",X"D8D1",X"D5D9",
      X"CDD0",X"CDC9",X"D6D4",X"D8D8",X"D0D4",X"CDCD",X"D2CD",X"DFDB",
      X"D6D8",X"D0D4",X"C6C9",X"CCC8",X"D6D1",X"D3D6",X"CDD0",X"CFC9",
      X"D6D4",X"D8D8",X"CED3",X"CCCC",X"D2CD",X"DFDB",X"CFD9",X"CDCB",
      X"CECE",X"DBD4",X"D3DA",X"CBCC",X"CAC4",X"D8D1",X"DBDC",X"5FA3",
      X"A05C",X"FEE4",X"F6FB",X"F2F3",X"F1F2",X"F1F1",X"F1F1",X"F4F1",
      X"F8F7",X"98D5",X"C49C",X"CACC",X"CAC9",X"CCC9",X"DECF",X"67CF",
      X"2C23",X"282B",X"2929",X"1E2A",X"8922",X"8C8F",X"8C8C",X"918F",
      X"9394",X"CDA4",X"D6D8",X"D0D4",X"C6C9",X"CCC8",X"D6D1",X"D3D6",
      X"CDD0",X"CFC9",X"D6D4",X"D8D8",X"CED3",X"CCCC",X"D2CD",X"DFDB",
      X"D8DA",X"D2D5",X"C9CD",X"D1CC",X"DAD6",X"D4D7",X"CDD1",X"D2CD",
      X"DBD8",X"DCDE",X"D3D8",X"CECF",X"D7D3",X"E0DE",X"D2DA",X"D2D0",
      X"D4D4",X"DDD8",X"D6DB",X"CED0",X"CDCD",X"BCCC",X"83AA",X"9B88",
      X"529A",X"9C4F",X"FAE1",X"F4FA",X"F2F4",X"F1F1",X"F0F1",X"F8F3",
      X"B9F1",X"AC8E",X"CAC8",X"CACA",X"CAC9",X"CCC9",X"D5D6",X"2378",
      X"2925",X"2628",X"2927",X"2B29",X"2422",X"986E",X"918F",X"9393",
      X"9394",X"9692",X"D8BF",X"D2D5",X"C9CD",X"D1CC",X"DAD6",X"D4D7",
      X"CDD1",X"D2CD",X"DBD8",X"DCDE",X"D3D8",X"CECF",X"D7D3",X"E0DE",
      X"DADB",X"D8D9",X"CED2",X"D8D2",X"DFDC",X"D6DC",X"D2D5",X"D6D1",
      X"E0DD",X"E1E2",X"D7DC",X"D1D3",X"DCD9",X"E0E0",X"D9DD",X"D7D7",
      X"DCD8",X"D6DB",X"B7C2",X"90AB",X"7C86",X"9483",X"C4A8",X"E0D5",
      X"41B9",X"1E16",X"A259",X"F7DA",X"F6FA",X"F1F2",X"F4F1",X"E2FA",
      X"96A4",X"D3BB",X"C9CC",X"C8C9",X"CBCA",X"D5CC",X"89D8",X"2325",
      X"2626",X"2726",X"2A2A",X"2A2A",X"262D",X"775A",X"9A84",X"9596",
      X"9494",X"9595",X"A193",X"D8C4",X"CED2",X"D8D2",X"DFDC",X"D6DC",
      X"D2D5",X"D6D1",X"E0DD",X"E1E2",X"D7DC",X"D1D3",X"DCD9",X"E0E0",
      X"DEE0",X"DCDC",X"D2D6",X"DBD7",X"E3E0",X"DCE0",X"D6DA",X"D9D6",
      X"E2DF",X"E2E3",X"D9DE",X"D1D7",X"D6D3",X"DADA",X"DCDB",X"D2D9",
      X"95B6",X"A69C",X"A5A9",X"A6A1",X"BEB0",X"DBD0",X"CBD7",X"AFC0",
      X"2361",X"272C",X"742B",X"9D85",X"F9DB",X"F5FA",X"F5F7",X"93C7",
      X"C8A0",X"CED2",X"CBCA",X"C9C8",X"CECC",X"D0D5",X"368E",X"2927",
      X"2627",X"2726",X"2A2A",X"2927",X"2B32",X"DB68",X"7DAD",X"9B8B",
      X"9695",X"9C9A",X"9595",X"A696",X"D2C0",X"DBD7",X"E3E0",X"DCE0",
      X"D6DA",X"D9D6",X"E2DF",X"E2E3",X"D9DE",X"D5D7",X"E0DD",X"E0E3",
      X"E0E1",X"DCDF",X"D4D8",X"DDD6",X"E5E3",X"DFE3",X"D9DC",X"D9D7",
      X"E1DF",X"E1E3",X"CAD7",X"91A8",X"978E",X"9997",X"A09C",X"6789",
      X"EAAF",X"F7FB",X"E2E4",X"E3E0",X"DBE3",X"ADCB",X"788E",X"967B",
      X"2357",X"2B30",X"8C25",X"86B5",X"9876",X"EDD6",X"A2DA",X"A987",
      X"D0D0",X"CDCD",X"CCCD",X"CCCC",X"DAD1",X"73C2",X"2E2E",X"262D",
      X"2626",X"2A29",X"292B",X"2927",X"3437",X"D32F",X"F2FF",X"7BAE",
      X"987A",X"9898",X"9797",X"9797",X"9B94",X"DDB9",X"E5E3",X"DFE3",
      X"D9DC",X"D9D7",X"E1DF",X"E1E3",X"DBDE",X"D8D9",X"E2DF",X"E0E2",
      X"DFE0",X"D9DE",X"CED2",X"D9D2",X"E3DC",X"DBE1",X"D6D9",X"D7D4",
      X"DFE0",X"B0DF",X"D38E",X"F2EE",X"F6F3",X"F0F6",X"E3F2",X"B29B",
      X"FFFF",X"D2ED",X"B4C0",X"9FA8",X"8696",X"7B7A",X"AE93",X"D2C4",
      X"1D6A",X"2B2B",X"7520",X"CDD0",X"84AE",X"9380",X"9286",X"D1BD",
      X"CECE",X"CBCB",X"CBCE",X"D4CD",X"B8DA",X"2363",X"322B",X"332F",
      X"2828",X"2C2C",X"282B",X"3128",X"3A3C",X"8B26",X"FFFA",X"EDFF",
      X"77B5",X"8B7A",X"9695",X"9596",X"8D91",X"A08E",X"E1C6",X"DBE1",
      X"D6D9",X"D7D4",X"DFE0",X"DFDF",X"D6DC",X"D5D4",X"E0DB",X"E1E2",
      X"DBDC",X"D4D9",X"C8CC",X"D1CC",X"E0DB",X"D7DF",X"D2D4",X"D1D0",
      X"DCDA",X"7896",X"FFEF",X"FFFF",X"FFFF",X"FFFF",X"BBFF",X"B67E",
      X"97B1",X"717C",X"7471",X"7771",X"9883",X"CCB5",X"D8D7",X"DFD6",
      X"1A73",X"2427",X"701F",X"D4C8",X"CFD6",X"B3BD",X"D0BE",X"CDD1",
      X"CDCD",X"CCCD",X"CDCC",X"D1D5",X"4E9B",X"2F27",X"7531",X"B7A9",
      X"2C89",X"2C2B",X"292A",X"3D31",X"3C3E",X"612C",X"DD9E",X"FFFF",
      X"F6FF",X"6DB7",X"9051",X"9299",X"8A8D",X"8F8B",X"9896",X"CCB0",
      X"D2D4",X"D1D0",X"DCDA",X"E0E0",X"D3DA",X"CFCE",X"DAD5",X"E1E0",
      X"D6D4",X"CCD4",X"C5C6",X"CCC8",X"DBD5",X"D3D8",X"CCCF",X"CCCB",
      X"8ED3",X"F56A",X"FEFF",X"FBFC",X"FCFB",X"FFFC",X"6ACD",X"B28B",
      X"ACB1",X"B9AB",X"CBC0",X"CFCF",X"D5D2",X"D1D3",X"CFD0",X"E0D1",
      X"1973",X"2326",X"6115",X"D4CD",X"CDCD",X"D6D3",X"CFD2",X"CDCC",
      X"CFCD",X"CECE",X"D8CE",X"74C2",X"242A",X"3435",X"B451",X"CEC3",
      X"6CC4",X"2924",X"3129",X"3E3B",X"3C3E",X"A62E",X"93BC",X"FDC3",
      X"FFFF",X"F4FF",X"85B8",X"836F",X"898A",X"8B8A",X"9591",X"9093",
      X"BBA0",X"CCCB",X"D8D3",X"DBDF",X"CED4",X"CDCC",X"D5D0",X"DFDB",
      X"D2CF",X"C9D1",X"C4C3",X"CDCA",X"D5CE",X"CFD4",X"C9CC",X"CCC8",
      X"559F",X"FFE8",X"FBFD",X"FBF9",X"F8F9",X"F0FF",X"B78D",X"FEFB",
      X"E4FB",X"D4D8",X"D3D3",X"D1D1",X"CDCE",X"CDCB",X"CECE",X"E7D4",
      X"1C7C",X"2824",X"2A1A",X"D9AF",X"CACD",X"D1CE",X"CDD1",X"CECD",
      X"D0CE",X"D5D1",X"A5D7",X"1952",X"251D",X"312C",X"AD68",X"C4A0",
      X"81CD",X"2B1F",X"3B31",X"3F3F",X"383F",X"D435",X"DEFF",X"A79D",
      X"FFE1",X"FFFF",X"FEFF",X"A0DA",X"7573",X"9086",X"908E",X"8D8F",
      X"8C8E",X"AE94",X"D5C6",X"D6DB",X"CCCD",X"D0CD",X"D1CF",X"DBD6",
      X"D5D8",X"D4D4",X"D5D5",X"D2D2",X"DFD5",X"D3DE",X"CACC",X"BCCB",
      X"D342",X"FEFF",X"FCFB",X"F9F9",X"FBF8",X"C2FF",X"FAA9",X"FCFE",
      X"D6F3",X"CACC",X"C9CA",X"CCCB",X"CECD",X"CACC",X"CECC",X"E4D2",
      X"1F86",X"2B27",X"1227",X"D169",X"CDD7",X"CFCD",X"CECE",X"CDCD",
      X"D3CF",X"CFDE",X"2F87",X"2117",X"2728",X"4822",X"9A7C",X"A797",
      X"7DB8",X"3426",X"403D",X"4041",X"3440",X"EF4D",X"FFFF",X"B4F6",
      X"C493",X"FFF4",X"FFFF",X"FFFF",X"B1EF",X"5D6C",X"947F",X"9096",
      X"8D8D",X"8F8D",X"AC91",X"DED0",X"D0D4",X"CBCE",X"D9D2",X"E1E1",
      X"D6DA",X"CDD2",X"CDCD",X"CECE",X"DAD2",X"CFD7",X"CDCC",X"5ACC",
      X"FFBC",X"FAFF",X"F9FB",X"F9FB",X"FFFC",X"A8EC",X"FEE1",X"F9F8",
      X"DDF8",X"CDCB",X"CBCD",X"CECA",X"CDCE",X"CDCB",X"D0CE",X"E7D2",
      X"2193",X"2C2A",X"212B",X"961F",X"D3DE",X"CECE",X"CFCE",X"CDCC",
      X"D8D4",X"61AD",X"1F22",X"2428",X"2C29",X"934F",X"C7C3",X"C3C6",
      X"61A2",X"3A2E",X"4240",X"4042",X"2E3E",X"FF6B",X"FEFF",X"FEFE",
      X"A5D8",X"C3AA",X"FBE3",X"FFFF",X"FFFF",X"BEF8",X"4F76",X"9576",
      X"8F8D",X"8E8F",X"938E",X"9D95",X"CFB5",X"CFCF",X"D3CF",X"DBD9",
      X"D9DE",X"CBD2",X"C9C8",X"CECB",X"D6D3",X"CED4",X"D0CD",X"9F93",
      X"FFFF",X"FBFD",X"FBFB",X"FBF9",X"FFFE",X"B7C3",X"FCFE",X"F8F7",
      X"E9FA",X"CCCD",X"CCCD",X"CBCB",X"CBCB",X"CCCA",X"D1D0",X"E4D3",
      X"1F88",X"2A28",X"2D2C",X"4612",X"DBBB",X"CECE",X"CED0",X"DBD4",
      X"85C8",X"1B37",X"2D29",X"202E",X"6429",X"9164",X"CCC8",X"CECB",
      X"82C8",X"4A5D",X"423D",X"3F40",X"2D3C",X"FFA5",X"FDFE",X"FDFB",
      X"F7FF",X"BBD8",X"AEA7",X"F2CE",X"FFFF",X"FFFF",X"D4FE",X"578B",
      X"977A",X"8D8E",X"918E",X"8E91",X"978C",X"CEC2",X"D2CE",X"D9D6",
      X"DBDF",X"CFD6",X"CCCC",X"D1CE",X"DAD7",X"D1D6",X"BCD2",X"EB6E",
      X"FFFF",X"F9FB",X"FBFC",X"FAF9",X"EFFF",X"DEA5",X"F9FE",X"F8F6",
      X"F5FA",X"CBD9",X"CDCF",X"CACB",X"CBCA",X"CECC",X"D1CF",X"E4D7",
      X"1C74",X"2A26",X"2C2C",X"1722",X"D271",X"CED6",X"D7D0",X"A4D5",
      X"2158",X"2D20",X"2A2A",X"1C2A",X"A072",X"6258",X"C9C3",X"CBB9",
      X"BED4",X"ABBB",X"3E36",X"3F3F",X"3638",X"FFD9",X"FCFC",X"F7FA",
      X"FEF9",X"FCFF",X"CFE9",X"B0B1",X"E2C4",X"FEFB",X"FFFF",X"DDFF",
      X"7386",X"8E8D",X"9392",X"9293",X"8D8E",X"C790",X"D8D1",X"DDDF",
      X"DBDB",X"D5D9",X"D1D2",X"D6D4",X"DFD9",X"D8DE",X"69D2",X"DE8E",
      X"FDFF",X"FBFC",X"F9FC",X"FBF8",X"CFFF",X"FEB8",X"F8FA",X"F8F8",
      X"FBFA",X"D4EC",X"CECD",X"CCCD",X"CDCD",X"CFCD",X"D1CE",X"E4DB",
      X"1E69",X"2A27",X"2B2A",X"1F2C",X"9923",X"DADE",X"BFDE",X"2578",
      X"2816",X"242B",X"2A26",X"5024",X"C5BF",X"72A8",X"CAAC",X"C9B3",
      X"D3D7",X"CBDA",X"394A",X"3E3E",X"6133",X"FFFB",X"FCFB",X"F9FA",
      X"F9F9",X"FBFA",X"FEFC",X"DDFA",X"AABC",X"DABB",X"FEF4",X"FFFE",
      X"6FC7",X"9992",X"9696",X"9696",X"8F93",X"9E8C",X"DFC3",X"E2E4",
      X"D9D7",X"D8D9",X"D3D6",X"D7D5",X"E0D9",X"DDE1",X"918B",X"E7A3",
      X"FAFF",X"F9F9",X"F9FB",X"FDF8",X"B4F7",X"FEDA",X"F7F8",X"F8F8",
      X"FBF8",X"E3F8",X"CBCF",X"CCCE",X"CBCE",X"CFCE",X"D3D1",X"D6DE",
      X"1E4F",X"2928",X"2B2A",X"302F",X"5325",X"D2B6",X"51A0",X"211C",
      X"292D",X"6B29",X"B2A6",X"9A7E",X"CACC",X"BCCA",X"D0AD",X"D4D6",
      X"D1D9",X"DBD1",X"3199",X"393E",X"AD2F",X"FFFF",X"FCFC",X"F9FC",
      X"F8F9",X"F8F9",X"FAF8",X"FEFD",X"ECFC",X"BCD1",X"C4B2",X"F0E7",
      X"BDA9",X"B7DA",X"999F",X"9697",X"9294",X"9291",X"A296",X"DCBA",
      X"D9D7",X"D8D9",X"D2D4",X"D9D5",X"DFD9",X"D4E0",X"CC7C",X"FBA7",
      X"FBFF",X"FBFB",X"F7F9",X"FFF7",X"B0E4",X"FBF1",X"F6F7",X"F8F6",
      X"FAF8",X"F4FC",X"CADB",X"CCCC",X"CBCB",X"CECC",X"D6D0",X"B3E3",
      X"2231",X"2A29",X"2A2B",X"2425",X"2A24",X"5B50",X"2230",X"2924",
      X"242E",X"B94F",X"C6C8",X"BC9F",X"C7CA",X"CFCA",X"C8D0",X"DACB",
      X"BBDD",X"DB95",X"35C3",X"333D",X"F14C",X"FDFF",X"FBFC",X"F9FB",
      X"F9F8",X"F8F8",X"F8F8",X"F9F8",X"FCFA",X"FBFE",X"C0E2",X"D0C1",
      X"ECA5",X"FFFF",X"D1EF",X"A3B3",X"9497",X"9592",X"9996",X"9999",
      X"DBD9",X"D8DB",X"D2D4",X"D9D7",X"DFDC",X"C0DF",X"C6C1",X"FFB3",
      X"FBFE",X"FBFD",X"F9FA",X"FFF8",X"C2C2",X"F8FC",X"F8F7",X"F8F8",
      X"F9F8",X"FCFB",X"D3EE",X"CDCA",X"CCCD",X"CFCD",X"D7CF",X"87E7",
      X"2922",X"2B2B",X"272C",X"2020",X"2522",X"2124",X"2A29",X"2427",
      X"222D",X"C779",X"ADC1",X"C28E",X"B9CA",X"D6C6",X"99D4",X"D490",
      X"CCE1",X"DAAC",X"3BCB",X"2F3A",X"FFA1",X"FBFF",X"FBFC",X"FAFB",
      X"F9F8",X"F8F8",X"F8F8",X"F8F8",X"F7F8",X"FBF9",X"FCFE",X"C9F5",
      X"FBA4",X"FCFE",X"FFFD",X"F2FD",X"BBDB",X"9699",X"9995",X"999C",
      X"DCDD",X"D3D8",X"CCCD",X"D5D0",X"E0DC",X"A1DE",X"B0F0",X"FFD0",
      X"FCFD",X"FBFB",X"F9F8",X"F4FD",X"D7A3",X"F6FE",X"F8F7",X"F6F7",
      X"F8F8",X"FBF8",X"ECFB",X"CAD1",X"CECC",X"D5CF",X"D9D0",X"64E0",
      X"2A22",X"2827",X"232A",X"2522",X"2526",X"2726",X"2C2B",X"2827",
      X"1E29",X"CB7A",X"C2CD",X"C696",X"C5CF",X"DAC9",X"BAD8",X"CD84",
      X"D1E1",X"DAC1",X"2FAD",X"5038",X"FFEB",X"FCFD",X"FBFB",X"FAFA",
      X"F9F8",X"F8F9",X"F8F8",X"FAF8",X"F9FA",X"F8F8",X"FBF8",X"B6FF",
      X"FFB2",X"FBFD",X"F9F9",X"FFFD",X"FEFF",X"C7E7",X"9BA7",X"999C",
      X"D9DD",X"CAD2",X"C4C6",X"C9C7",X"DFD8",X"9FD0",X"A8FD",X"FFE0",
      X"F9FC",X"F9FB",X"F8F9",X"DCFF",X"EDA0",X"F7FB",X"F8F8",X"F8F8",
      X"F8F8",X"F9F8",X"F9FA",X"D1E9",X"CFCC",X"D4D1",X"DAD2",X"47CC",
      X"2921",X"2B2B",X"302A",X"2127",X"2924",X"2528",X"2324",X"2A23",
      X"212E",X"C567",X"BCCD",X"C587",X"D6D2",X"D7D3",X"DAD9",X"AFBB",
      X"C9DB",X"D4C6",X"355E",X"9230",X"FFFF",X"FBFC",X"FBFC",X"FAFA",
      X"FAFA",X"F8F9",X"F9FA",X"F9F8",X"F9FA",X"F8F8",X"FEF8",X"A3F9",
      X"FFDC",X"F9FB",X"F9FB",X"F8F9",X"FDFB",X"FFFF",X"D7F5",X"9FBA",
      X"D5DA",X"C8CF",X"C5C5",X"C9C8",X"DED5",X"C593",X"A6F5",X"FFEF",
      X"FBFB",X"F9FB",X"F9F9",X"BFFF",X"FDB3",X"F8F9",X"F9F8",X"F7F8",
      X"F8F8",X"F9F8",X"FAF8",X"E6F9",X"CED1",X"D1CF",X"DFD2",X"34B4",
      X"2B23",X"272B",X"6F35",X"1F36",X"2B2C",X"2526",X"2122",X"2523",
      X"292E",X"863F",X"9BBA",X"A363",X"D6CE",X"D9D6",X"DED9",X"A0D3",
      X"B0B8",X"C0D1",X"3228",X"E446",X"FEFF",X"FBFC",X"FBFA",X"F8F9",
      X"F9F9",X"F8F8",X"F9F9",X"F9F8",X"F9FA",X"F8FA",X"FFFB",X"A4DA",
      X"FFF7",X"F9F9",X"FBFB",X"FBFB",X"F8F9",X"FCFB",X"FFFE",X"DDFD",
      X"D6D8",X"CDD2",X"CAC9",X"D0CD",X"D2D8",X"E95F",X"B8ED",X"FEFD",
      X"FBFB",X"F9FB",X"FDF9",X"A3F9",X"FFC9",X"F8F9",X"F9F9",X"F8F9",
      X"F7F8",X"F7F6",X"F8F8",X"FAFB",X"D0E4",X"CDCF",X"E3D2",X"2BA1",
      X"2C27",X"1E2A",X"B85F",X"2037",X"2A2F",X"2625",X"2626",X"2727",
      X"2526",X"2620",X"2A35",X"891E",X"D8CD",X"CDD7",X"D4CE",X"ACD4",
      X"C376",X"74D8",X"2E28",X"FF96",X"FCFE",X"FBFB",X"FAFC",X"FCFA",
      X"FAFA",X"F9F8",X"F8F8",X"FAF9",X"F9FA",X"F8F8",X"FFFB",X"BEBF",
      X"FEFF",X"FBFB",X"FCFB",X"F9FC",X"F9F9",X"FAF9",X"FAF8",X"FEFC",
      X"D9D8",X"D5DA",X"CCCF",X"D5D0",X"B7DE",X"FF61",X"C4EB",X"FEFE",
      X"F9FB",X"F8FA",X"FFF8",X"96E4",X"FEE5",X"F9FA",X"F9F9",X"FAFA",
      X"F7F8",X"F7F6",X"F8F8",X"FBF9",X"E1F9",X"CED0",X"E2D0",X"2586",
      X"2D2A",X"2523",X"C8AD",X"1C2F",X"282E",X"2929",X"2828",X"2627",
      X"2A25",X"2B29",X"393A",X"A52F",X"DAD7",X"AFD9",X"B59D",X"A2AF",
      X"E0BC",X"2DB8",X"532C",X"FFEB",X"FCFD",X"FAFA",X"FAFA",X"FBFA",
      X"FAFB",X"F9FA",X"FAFA",X"F8F8",X"F9F9",X"F8F8",X"F8FC",X"D8AB",
      X"FDFF",X"FBF9",X"FDFA",X"FBFC",X"F9FA",X"FBF9",X"F8F9",X"F9F9",
      X"DDD9",X"DDE1",X"D5D7",X"DED9",X"ABDF",X"FF84",X"D0E6",X"FEFE",
      X"FBFB",X"F7FA",X"FFF8",X"A1C0",X"FCFB",X"F9F9",X"F9F9",X"FAF9",
      X"F8F9",X"F8F8",X"F8F9",X"FAF8",X"F7FD",X"D0E1",X"DFD1",X"2576",
      X"2928",X"611B",X"C3EB",X"1931",X"2827",X"2729",X"2926",X"292B",
      X"262A",X"552F",X"323D",X"D048",X"D9DC",X"D2D8",X"D1D1",X"D3CC",
      X"CEE4",X"2B4B",X"BE38",X"FEFF",X"FCFC",X"F9FA",X"FAFA",X"FAFB",
      X"FBFA",X"FBFB",X"FAFA",X"F8FA",X"F9F8",X"F8F9",X"E8FE",X"EBA0",
      X"FCFF",X"F9F9",X"FAF9",X"FBFB",X"FBFB",X"FBFB",X"FAFB",X"FBFA",
      X"DDDA",X"DFE0",X"DAD9",X"E3DE",X"6FDE",X"FFB4",X"D8E3",X"FEFE",
      X"FBFB",X"F7FA",X"FFFD",X"B89B",X"FBFE",X"F9FB",X"F9F9",X"FAF9",
      X"F8FA",X"F8F8",X"F8F8",X"FAF9",X"FDFC",X"E1F7",X"D4D3",X"225E",
      X"1D29",X"B335",X"BBED",X"1831",X"2424",X"2524",X"2B27",X"3030",
      X"1C2B",X"CD4E",X"2864",X"9A40",X"DACE",X"D9D8",X"DCDA",X"E2DF",
      X"62CD",X"2A2E",X"FF81",X"FBFF",X"FBFC",X"FAFA",X"F9F8",X"FBFB",
      X"FAFB",X"FAFA",X"FAF8",X"FAFB",X"F8FA",X"F9F8",X"C5FF",X"FFA2",
      X"F9FD",X"FBFB",X"FBFB",X"FBFC",X"F9FB",X"FBFB",X"FAF9",X"FFFE",
      X"DDDC",X"DADD",X"D6D6",X"DCD8",X"64DF",X"FFD2",X"D0DB",X"FCFF",
      X"F9FA",X"F8FA",X"E6FF",X"DF86",X"FAFE",X"F9F9",X"F9F9",X"F8F9",
      X"F8F8",X"F8F8",X"FAF9",X"F9FA",X"FCFA",X"F8FC",X"CCE6",X"2151",
      X"3423",X"DB92",X"A8E3",X"1D25",X"2222",X"2827",X"2F2A",X"3334",
      X"1A2B",X"FF88",X"40D8",X"2B2A",X"DAB4",X"D8DB",X"DDDA",X"BFD4",
      X"3050",X"5D2D",X"FFF1",X"FBFD",X"FAFB",X"FAFA",X"FAF9",X"FAFA",
      X"FAFA",X"F8F9",X"FAF8",X"FAFA",X"F9FA",X"FCF8",X"A7FE",X"FFB9",
      X"F9FD",X"FBFB",X"FBFB",X"F9FB",X"F9F9",X"F9FB",X"FFF8",X"E0FF",
      X"DADC",X"D6D9",X"CED1",X"D4D0",X"55C3",X"FFEC",X"C1DC",X"FEFF",
      X"FBF8",X"FAFA",X"C6FF",X"FB92",X"F8FC",X"F9F9",X"F9F9",X"F8F9",
      X"F8F8",X"F8F8",X"FAFA",X"F9FA",X"FBF8",X"FEFB",X"D3FD",X"2149",
      X"8226",X"D1D8",X"9EE0",X"1E22",X"2A25",X"2D2F",X"322D",X"3232",
      X"2F24",X"FFCD",X"A9FF",X"3230",X"A13B",X"D4C3",X"B2CD",X"3D7D",
      X"3232",X"CC35",X"FEFF",X"FBFB",X"FAFB",X"FAFA",X"F8F8",X"FAF9",
      X"FAFA",X"FAFA",X"FAFA",X"F9FA",X"FAFA",X"FEF8",X"94ED",X"FFDC",
      X"FBFC",X"FBFA",X"FBF9",X"F8FB",X"FBF9",X"FBFB",X"FFFE",X"BBDC",
      X"D7D9",X"D2D4",X"CBCE",X"D1CD",X"66C1",X"FFFE",X"BADE",X"FFFB",
      X"FBF9",X"FCFA",X"B1FF",X"FFAD",X"F8F9",X"F8F8",X"F8F9",X"F8F8",
      X"FAF8",X"F9FA",X"FAFA",X"F9FA",X"FAF9",X"FDFA",X"D9FF",X"2044",
      X"D069",X"CED1",X"98E9",X"251F",X"2E2A",X"2B2E",X"312D",X"3132",
      X"6E18",X"FFFF",X"FEFF",X"3273",X"2F36",X"7F4C",X"3263",X"3831",
      X"2D37",X"FF8C",X"FCFF",X"FBFB",X"FAFA",X"F9FA",X"F8F8",X"F9F9",
      X"FAF8",X"FAFA",X"FAFA",X"F9F9",X"F8F9",X"FFF9",X"98D8",X"FFF4",
      X"FBF9",X"FCF9",X"F9FB",X"F9F9",X"FAFA",X"FBF8",X"E9FF",X"E7B5",
      X"D6DA",X"D0D2",X"CBCC",X"D0CC",X"7CAC",X"FFFF",X"ACE0",X"FFF8",
      X"FBFB",X"FEF9",X"98FD",X"FFC8",X"F8FA",X"F8F8",X"F8F8",X"F8F8",
      X"F8F8",X"F9F9",X"FAFA",X"FAFB",X"F8F8",X"FBF8",X"D4FF",X"5235",
      X"DCCC",X"E7D6",X"A1FF",X"2B22",X"2E2A",X"282F",X"2E28",X"2731",
      X"BE23",X"FEFF",X"FFFE",X"49E0",X"3E35",X"3539",X"3C38",X"3C3F",
      X"652E",X"FFF8",X"FBFD",X"FAFA",X"FAFA",X"F9FA",X"F8F8",X"F9F9",
      X"F9F8",X"FAFA",X"FAFA",X"F9FA",X"F9F9",X"FFFC",X"AFC0",X"FDFF",
      X"F9F9",X"FCF9",X"F9FB",X"F9F8",X"F8FB",X"FDF8",X"BCFB",X"FFC8",
      X"D7DC",X"CFD3",X"C9CB",X"CFCB",X"94AE",X"FFFF",X"A7E0",X"FFF2",
      X"F7F9",X"FFFB",X"84E9",X"FFDE",X"F9F9",X"F8F8",X"F8F8",X"F8F8",
      X"F8F8",X"F9F9",X"FAF9",X"FAFB",X"FAFA",X"FCFA",X"BAFF",X"AE2E",
      X"F5FE",X"FFFB",X"A4FF",X"2B26",X"2E2E",X"2B2D",X"2E26",X"162A",
      X"FB70",X"FEFF",X"FFFD",X"ABFF",X"3836",X"3F3E",X"3D3E",X"313E",
      X"D747",X"FDFF",X"FAFA",X"FAFA",X"FAFA",X"FAFA",X"F9FA",X"F9F9",
      X"F9F9",X"FAFA",X"FAFA",X"FAFA",X"F8F8",X"FDFE",X"CEA6",X"FAFF",
      X"F9F9",X"F9F9",X"F9FB",X"FAF8",X"F9FB",X"FFFB",X"B1DC",X"FFF4",
      X"D6DA",X"D0D3",X"CCCE",X"D4CF",X"A8B5",X"FFFF",X"A2EB",X"FFEB",
      X"F9F9",X"FFF9",X"83D0",X"FEF3",X"F8F7",X"F8F8",X"F8F8",X"F8F8",
      X"F9F8",X"F9F9",X"F9F9",X"FAFB",X"FAFA",X"FDFA",X"C8FF",X"D958",
      X"FFFF",X"FFFF",X"A3FF",X"2A26",X"2E30",X"2B2F",X"2B2A",X"371F",
      X"FFD1",X"FCFF",X"FEFD",X"FEFF",X"3083",X"3E39",X"3F3F",X"3038",
      X"FFAD",X"FBFF",X"FCFB",X"FAFA",X"F9F9",X"FAFA",X"FAFA",X"F9F9",
      X"F8FA",X"FAF8",X"FAFA",X"FAFA",X"F8F8",X"E5FF",X"E994",X"FAFF",
      X"FBF9",X"F9FB",X"FBFB",X"F9FB",X"FBF9",X"F7FD",X"D5B7",X"FBFF",
      X"D9DC",X"D8D8",X"D5D5",X"DFDA",X"C0BB",X"FFFF",X"9AF5",X"FFDF",
      X"F9FB",X"FFF9",X"98BC",X"FBFD",X"F8F6",X"F8F9",X"F8F8",X"F7F8",
      X"F8F8",X"F9F8",X"F9FA",X"F9FA",X"FAF8",X"FBFA",X"E2FF",X"E688",
      X"FEFF",X"FFFE",X"AAFF",X"2424",X"2B2B",X"2A2B",X"2A2B",X"8C1C",
      X"FFFF",X"FDFF",X"FFFC",X"FFFE",X"5CF3",X"3B2D",X"4041",X"752E",
      X"FFFF",X"FAFD",X"FBFB",X"FAFB",X"F9F9",X"FAFA",X"FAF9",X"FAFA",
      X"FAFA",X"FAF8",X"FAFA",X"FAFA",X"FAF8",X"C4FF",X"FC9A",X"FBFF",
      X"FBFB",X"FCFA",X"FBFB",X"F9F9",X"FCF9",X"D5FF",X"F8B2",X"FBFD",
      X"DDDD",X"DCDE",X"D9DA",X"E5DE",X"D7BF",X"FFFF",X"9DFC",X"FFD0",
      X"FBFA",X"FFFE",X"AEA3",X"FAFF",X"F8F8",X"F8F9",X"F8F8",X"F8F8",
      X"F9F9",X"F9F9",X"FAFA",X"F8F9",X"FBF8",X"F8F9",X"D4FF",X"F594",
      X"FEFF",X"FFFE",X"BCFF",X"202B",X"2A26",X"292A",X"1E27",X"DE40",
      X"FFFF",X"FEFD",X"FDFD",X"FEFD",X"E0FF",X"3045",X"373F",X"DF3D",
      X"FEFF",X"FCFB",X"FBFA",X"FAFB",X"FAFA",X"F8F8",X"FAF8",X"FBFB",
      X"FAFA",X"F7F8",X"FAF9",X"FAFB",X"FBF9",X"B1FF",X"FFAD",X"FCFF",
      X"F9F9",X"FBFC",X"F9FB",X"F8FA",X"FEF8",X"B1FB",X"FFD0",X"F9FB",
      X"DBDA",X"DBDD",X"D3D6",X"DFD7",X"E1BA",X"FFFF",X"A5FF",X"FFC4",
      X"FAF9",X"F8FF",X"CE92",X"F9FF",X"FAFA",X"F8FA",X"F8F8",X"F9F9",
      X"F9F8",X"F9F9",X"F8F9",X"F8F8",X"F8F8",X"FAF8",X"C2FF",X"FFA2",
      X"FEFF",X"FFFF",X"A1FF",X"2627",X"292C",X"2529",X"2720",X"FFAE",
      X"FFFF",X"FBFC",X"FCFC",X"FDFD",X"FFFF",X"44CD",X"3234",X"FF97",
      X"FEFF",X"FAFC",X"FAFA",X"FAF9",X"FBFA",X"F8FB",X"FAF9",X"FCFB",
      X"FBFB",X"FAFB",X"FBFA",X"FAFB",X"FEFA",X"A2FE",X"FFC1",X"FDFE",
      X"FCFD",X"FDFA",X"FBFA",X"F8F9",X"FFFB",X"A5D8",X"FEF4",X"FAF8",
      X"D9DE",X"D3D6",X"CCCD",X"D8D2",X"EB9D",X"FEFF",X"ADFF",X"FFB4",
      X"F9F8",X"E8FF",X"E490",X"F7FF",X"FAF8",X"F9F9",X"F8F8",X"F9F9",
      X"F9F9",X"F9F9",X"F8F9",X"F8F8",X"F8F8",X"FAF8",X"B7FE",X"FFBF",
      X"FDFF",X"FFFF",X"46DC",X"2A1F",X"292B",X"262A",X"6719",X"FFFF",
      X"FDFD",X"FCFA",X"FDFC",X"FDFD",X"FFFE",X"90FF",X"6B2B",X"FFF9",
      X"FDFD",X"FAFB",X"FAFA",X"FAFA",X"FBFB",X"FAFB",X"FBFB",X"FBFA",
      X"FBFB",X"FBFB",X"FBFC",X"FAFA",X"FFFA",X"8FF1",X"FFDC",X"FCFE",
      X"FDFC",X"FDFD",X"FBFC",X"FCF7",X"FCFE",X"CEB0",X"FAFF",X"F9F9",
      X"D6D9",X"CED2",X"C5C8",X"D0CB",X"F08C",X"FEFF",X"BBFF",X"FFA4",
      X"F8FB",X"C9FF",X"F899",X"F8FD",X"F8F8",X"F9F9",X"F9F9",X"F9F9",
      X"F8F9",X"F9F8",X"F8FA",X"F8F8",X"F9F9",X"FBF8",X"A9FC",X"FFD6",
      X"FFFF",X"FEFF",X"176F",X"2826",X"2928",X"272D",X"A620",X"FFFF",
      X"FDFC",X"FBFB",X"FCFC",X"FBFC",X"FFFA",X"A4FD",X"EC9A",X"FEFF",
      X"FCFC",X"FAFB",X"FAFA",X"FBFA",X"FBFB",X"FAFB",X"FAFA",X"FBFA",
      X"FBFB",X"FBFB",X"FAFB",X"FAFA",X"FEF9",X"87D3",X"FFEF",X"FBFC",
      X"FCFD",X"FAFA",X"FBFC",X"FCF7",X"DEFF",X"F3A8",X"F8FF",X"FAF9",
      X"D6DA",X"CBD0",X"C2C4",X"C1C7",X"F581",X"FEFF",X"CEFF",X"FDA2",
      X"FCFE",X"ABFF",X"FFA7",X"F7FB",X"F8F8",X"F9F9",X"F9F9",X"F9F9",
      X"F8F9",X"F8F8",X"F9F8",X"F8F8",X"F9FA",X"FDF8",X"A1EE",X"FFE7",
      X"FFFF",X"ADFF",X"2120",X"2628",X"2A26",X"232C",X"BD24",X"FFFF",
      X"FDFD",X"FEFE",X"FDFE",X"FDFD",X"FFFE",X"B1D1",X"FFFC",X"FDFE",
      X"FCFC",X"FAFB",X"FCFA",X"FCFB",X"FAFB",X"FAF9",X"FAFA",X"FAFA",
      X"FBFA",X"FBFB",X"FAFB",X"FAF9",X"FFFC",X"9CBF",X"FFFA",X"FCFB",
      X"F9FC",X"FBFC",X"FBFC",X"FBF8",X"B6FE",X"FFC8",X"F9FB",X"FAFA",
      X"DADE",X"CFD5",X"C5C7",X"BFC9",X"FC86",X"FAFC",X"DDFC",X"EF97",
      X"F7FC",X"99F7",X"F8BE",X"F0F3",X"F1F1",X"F2F2",X"F1F2",X"F2F1",
      X"F2F2",X"F4F4",X"F2F2",X"F1F1",X"F2F2",X"F8F1",X"9DDD",X"F8EE",
      X"F9F8",X"52E7",X"311F",X"2F2D",X"3130",X"2830",X"B829",X"F9F9",
      X"F6F8",X"F8F7",X"F8F7",X"F7F7",X"ECF8",X"DDB1",X"F5F8",X"F5F5",
      X"F5F4",X"F3F5",X"F5F3",X"F4F4",X"F4F5",X"F2F2",X"F4F3",X"F4F4",
      X"F5F5",X"F5F5",X"F6F6",X"F4F4",X"F8F5",X"AFA7",X"F9F9",X"F4F4",
      X"F5F4",X"F6F6",X"F4F6",X"F9F3",X"ABD9",X"F9EC",X"F3F2",X"F4F5",
      others=>(others=>'0')
      );
  type state_type is(IDLE,WR1, WR2,WR3,WR4);
  constant offset : integer := 8;
  constant dlen : integer := 8192;
  signal state,state_next: state_type;
  signal ram_addr, ram_addr_next: unsigned(13 downto 0) ;
  signal read_mode : std_logic := '0';
begin
    process(clk)
	begin
      if reset = '1' then
        ram_addr <= (others=>'0');
        state <= IDLE;
        read_mode <= '0';
      elsif falling_edge(clk) then
        ram_addr<= ram_addr_next;
        state <= state_next;
        if finish = '1' then
          read_mode <= '1';
        else
          read_mode <= read_mode;
        end if;
        
      end if;
      
	end process ; -- 
    
    -- combinational circuit
    process(start, state, ram_addr, finish)
    begin
      state_next <= state;
      ram_addr_next <= ram_addr;
      adv <= '1';
      cs <= '1';
      rw <= '1';
      --ready <= '0';
      case state is
        when IDLE=>
          da <= (others=>'0');
          if start = '1'  then
            --adv <= '0';
            ram_addr_next <= (others=>'0');
            --state_next <= WR1;
          elsif(ram_addr < dlen) then
            adv <= '0';
            da<= std_logic_vector(("0"&ram_addr&"0") + offset);
            state_next <= WR1;
          elsif ram_addr = dlen then
            -- start the sobel calcul
            adv <= '0';
            da <= X"0004"; -- trigger the sobel
            state_next <= WR1;
          elsif finish = '1' then
            ram_addr_next <= (others=>'0');
          end if;

        when WR1=>
          state_next <= WR2;
          da <= ram(to_integer(ram_addr));
          cs <= '0';
          if read_mode = '0' then
            rw <= '0';
          end if;
          
        when WR2=>
          state_next <= WR3;
          cs <= '0';
          if read_mode = '0' then
            rw <= '0';
          end if;

        when WR3=>
          state_next <= WR4;
          cs <= '0';
          if read_mode = '0' then
            rw <= '0';
          end if;
        when WR4=>
          state_next <= IDLE;
          cs <= '0';
          if read_mode = '0' then
            rw <= '0';
          end if;
          ram_addr_next<= ram_addr + 1;
      end case;
      
    end process;
    
end architecture ; -- arch
