mrsang@LEs-MacBook-Pro.local.909